PK   �XX��$x�  �    cirkitFile.json͜mo�H�����������W��t�6��t�=�]lbYl�HJN:�oQrl��ԑu"k�;2�:�sU,W�O��~�V�fݻ�{�o���Z���mݷ�ã�rr�XͶ���}}w;��4��l?޹�Y��[��j;+�ie�.Klֺ$k�m2�l�t����LS[���������E��ꚧ�普y�k^蚗�敮�TY6C�=����n�k_�3�\�I�%�K�$�U�LۦNڪ��|j�e3�u�yweՊ�lEY��,\QV�(KW��+��e�Z�i��������������������������Re��������&�6ܭ?�>����d���zY���G�xC­��J~��',?a��`���V?a��g��Ntb�}#lߘ`��r�,��e�������L����OY�RV?-?a�	����/����/c�������L�����Y�rV?-?a�	�����;�`�+X�����',?8_/��կd�������L`=���+V���O�OX~��3�������MY�����',?�7ߕO�{#�}��(0E�)���g�:���&�����h�?%���#���(0E�)��zg�:��lʨ)
LQ`�&����;3[3j�S��	��}F����������h�%g�:��lӨ)
LQ`�&\�qF��^��f�����h��6g�:��l٨)
LQ`�&\�tF�þ��ƍ����h¥gg���n,�ݨ)
LQ`�&\ xF��ލ��5E�)
Lф�0��uz%��XKC/����`1��{7�n��(0E.I>��a���ލ����h�g�:��XػQS���M�<��^��{7j�S��	7I���wca�FMQ`�S4�V�3z�n,�ݨ)
LQ`�&�0tF��ލ��5E�)�W(>�)��u׶�4IK7M��˓i�IR�iմmQ�i�;��Oj~|��I�w�q�w�]��z��'0��I��N�<�X%EP2%GP
�DP*e�Tݮx����j`���|��_a
X�
����aa�X�*��l�1��b�T�e��2Ul�*�L[��-S�)S��*>k_{H��G��H	�B����isl�����JK|����(=is�A��G��H�{�qTP�#��yT"��QA�����[�qTPi�t��G�>2	�o��QA�!��N|T��s�~{>�
*���㨠�Ge��qTPi�t��G�>�6��㨠��0 G�>b��pTPi�t�����	f�{�yX�<�|�QxG" �9�l$�l$��I!�aI�1�,ط�Òzc��(�#��ޘm���aI�1�lޑ�Ho�<� xXRo�?�w$
��Ђ� ��s�F�	M��ƌ� _��%�Ƽ�QxG� �1;-H"�aI�1Gmޑ Ho�T2xXRo�W�w$���ւt��s�F�	w�֫`�Z���ÒKV0mޑHo�_xXRo�_�w$0қ[�6Ҋ����qk�FZ�6��vlU;4�Òzc��(�#!�ޘ��5�ޘ�6
�H\�7��<,�7母�;l��kAK��k���D`@zc�Z��Òzc��(�#a�ޘ��J�ޘ�6
�H��7�	<,�7母�;��}y���]ӧ�r<�<�sl���i�9V�~����ŝΡG�J��dJ��J��Tʔ�:�x���|��_a
X�
����aa�X�*�L[hf��2Ul�*�L[��-SŖ�b�Tq�Tqz���� �4�~�
��t$��F�H�c�O ��F��HG�9hTP�#�& ��F��HG�9hTP�#� ��F��HG�9hTP�#3< ��F��HG�9hTP�#�p ��F��HG�9hTP�#�I@8�
*���sШ��Ge�pT"	�QA���@8�
*���sШ��G! ��F��HG�9hT�9�L�0��%��'�w,��ћ��F��F2�8�l$�l��؟$�p����F��`��l�0��%�Ɯ�Qx��9�1�,��aI�1�lޱpFo�BC*pXRo�E�w,���3�
����F��`���0��%���Qx��9�1S-��aI�1_mޱpFo�ZC*pXRo�]�w,��Y���kaHK.Y���Qx��9�1-��aI�1mޱpFonA�H+�FZ�ƭIiQ�8�ڱU�D8K��k����s0zc�ZR�Òzc��(�c��ޘ��Tతޘ�6
�X8�7毅!8,�7母�;����kaHK��k����s0zc�ZR�Òzc��(�c��ޘ��Tతޘ�6
�X8G��p=�WwM�������v֬��~�h�\g����mfw˺q�l��������7o��ٕ.�:��6+����d��76�<���ti�ܥ�m�ҵi�uY�T��$O+��y�es��*zsy��������w�/N��7�5zj�<�|�b^�k���'77_*�w���}�ի6V}o�u����eI�A_�'��7���VЇ�K
>z����~��9E�����A�A�����ۛ�}���v��i��~�zL�z�y�u�7b���6�k����4�}�l�)������}�l_)�O��3��͗O[���Hі�hkR�E)ڪmY��.E[�V;2Z�Ш�D��D��D��D��D��D��D���T[�iP��ef=�P�Z��#oo�(��b$��(�p��ʬBT��(U���'T�U��,cN�U�T�����j���+Q1�W�����3J�#�U�b0aR�J!*�a�*�)F��8<D�`֪��BTV�(UTS��Nqx�����*
Q1X��TQM1)��!*�o��'D�`E�RE5�H\���<D�b��u&J�#QP�b�d�"���#J�#1Oc ^Nn2> `��,c�MZ-	G�tpOG�2�2ZFNJ2Z^�2����s��!��pt`��@%�����	���������%i���0(d���e,I�%`��!@  �%���,c!GZ-�'�-�f0�j	�=ax�h	�=0�X8�VK��	�y@@FK���YƂ��� �'��������
i�|�0Pd�|�e,0H�%��_��/�!����xh�'\r�K�a��}=�X��h	�>a��h	�>0�X��VK��	l@@FK���Y�z�Z�ON2Z��2����}�����}`��`�����ʀ���������h�|�00d�|�e,��Q8����������|��n���=�fظ~�����ɰ�g��;�ߙ���w�K�]���p����LN��\N��lN��|���-�{ha�vha�vha�vha���"�\&�t��˿�q��]0�'x�`���7� x���Y���n9\mx�����D������-V�z�\l���"�a��?�{7�,��_����˶h�n�9��$k�U�en�2��I��i�?d��_���76f��k|�7��ݛ��^�clT��bn�\o����;��_߹~�p�ƻ���� ���Ͷ_�~�lV����ᷗ����~��O��P���������]�a��ǝ\wC��_n\��b��/�����~ѻvr���5|W����C��8<��J����K���b�X�~xS��eZTWe��o��W�<�Ym�yfR_�I��4Im�<��?R�e���������\N����W��Q�r����_Ӥ_�|��}�tR���^�k�����E���:8>}:��������ǫ�׹y:'��������x1/��m����T��=8����ǫ��y:�������������z������^�����xvp���}�ڡ�<���������������d��6�o'�o'�vw��b�J��P�M�K�u�'�q�0�ɪ��|���r���?��m��}vu�U���t��A�k���ش�V.ϻ]����I�9��Ub
_�Y1��ە�Ԯ�Ӯ(ˢ�۽Z��o7Y;��N�U���t�&u��I^�鴝���=�ͫ���o�O�~��=1��v�l�K)��9?2�~tͪ�Jj�Ebe^�+��]�>���_o�s����<m�.����)�_�)� Y�W27ټ��|�\o���t]ứ�����1<�NM�k���-�x���_��U���i9�c�_�9_��������������R&��y��j��m6��|)�S�]v���T������7u�1�W{�'	���`'��Ѭ����2r��楛Os�ɺ�W�IS/���HQUum�S�&Va�F��������ܷ�癯��ʝm�<sG+�4�-�&3�i:���1�T��ל�2�~���o'�׋�b��w����޾]]\����.>����o.��/n]�./���~u��#�?���y��h�^�q�ՋU�ww�޺v��l�?��k��������d?z��0�y���cE��qy�Yl�޷����d"W��������������������W��
��[)��"/��p��]Ji�L�eU��_4e�W�O���C�_�i[$�L�i��f>u'��O�����t]x��p���}����ڧ�T�����
�@��k�3�6���vW3�����c=$�.�zR��#�����/9�n7)��d�Ӊ�>o����lV7����q���w��ǟ��I��|����c��3���s���ϑ��~�z�z94��!p�F�^������?~����<��O�̇����n�Xm_������N�g����/~�}h7���7��m����k�+�ǯ���Y�>�,?Պ���;��Y7���q�̴X.�����~�G_m�z6��r����S/�[�{�u�;ꛛϓ��PK   �XX��8��9 z /   images/07769342-c5fd-4eb7-a5a5-41db20f507eb.pngT\\��׎�j[�4[AY6D������b+��
"�@Dd�����(5D@YVT� �M�(�+#�a�,�! {}�!��_�S���3���������|���op8ܷ��ZF8��|������&��K�_Hg��__]��߿v=i��I=G��y�p����󄙧��%O�9w;�BQppv��p��N���>vDc;�G����O�P��Ĕu�|��vj�����m�w=�*24��o�R���惐w����)\�|�e�|���5�������/W��*���ϯ]��H;h�I��G���W�놮صr�(���?�ޒ�f����ok�5)h48!�~b��Gݘ�8?5L�>��ޡ�o��p,^����V��"T�-�X��;Ğ��QU�əc'�f^Mɍ"��-r���g�2��K����ٓ�9�S�ǔ:y�C���(b����Jb���zE�'"%ʤ�����	��/F��#��a��ҕ��1�x��3��=H�ކ�=�	�z�7�=���%4���<��g�[l@��[���;u���Z&#�g�g��wV���{�����$Cl�.���9�Of[�������j]�Xob�y��CF�b�f �~�)�'�"f"v��ҋ�,x7�=��Z�,��ԅOz�3[H#�´�B^�����#k\,-�C��x�7/�:j�:
��brc��H�,�1�c��T�l�G=+�(��BQ�y53���i���xӣްo�g�8�3��SF��T�h�͎a�x_����Q����[�c?��r��E���V�MO*�|4Z����#n|�Pd��ޫi�6�Q/YC<P��}���^�Ǟ�t�\�&���6���fɍ�Il�p�?^
�Jh[��klp�� �U\��>���3�o��zﱭc�S`hݤ$��A!M���������/���3p�.��F.�����qpSE��Byy����<zA�=��e3žk3�ß�e)	�$�wpՉI����9�M�C�ןM2&�軛�Y�g�J-;��n��6��0�4�)��a�ԱTȞ20p�T+R�7֐���0��r96�vsm��%�FR޳��9O��"kvn��_r0�vL������=Ց��m(��a�Pk�}uCCC$dt$`��\�t���JR�J͗������g���x���e�[�I,p������\:�BR(�FRb�r�"I	�{n�å�$n�Y ��/���/����c8���o���{��TD"�"%}��ɸ��Z� Kb��e��2.���,V�|���2��͈N߁�7°���GX�����e�9_�Q���c>�,F�J�D���ʼ�;�8�d�/�M��z�&���r��t�m�m�Y�����Sgi�����?>���u��Kw��6��|>|�G�CW�/��ٻ�C�[/n�E�`XѨ�h��s�k����.�~ž�.[P�m���Ȧ.�t�E���nnnO~�
>������;���=��#l�'�~����B��n���l����6�u'	�"��Q�z�63�u�lW��k֦6d�ni�|/ �è�c�'`���T�GR;�vMׂZTox\�ֱ�ǯ�Ʒ�#1�����E�&>��lbs�o���8�����[����=Gqf�;���(�<�Xra��6$\�{��4Vɻ��|�Bb�7�����_R�� ���_�VWWK�[YY]��h/Ύ�N��555�7�?}"�"֫N/LЯ�������J9sw��
̀��
�BA/��Y�h@�v`������Ԥ_I{.g���?��n��`%�����1�SO>��}$='''$�67	��~w�oA�ĿP8'��F}4:,u�˗n-���D+��$wG��kc��k�8�x�XE��c�uNcf;�S�Q�]Ҕ�l�L�v�Ǐ�;3z9�sKO��^9a�y��H�J��U�Rh�L���@J�q���_�j���O.�-��E.��+l�{���#"y4`����_�O6S�MJJJ�{g�����"���զp�mw{��}���w3��/�=:�
�8�޸w�^r����+�QF#�9��+���/��r�=�к.�;�~�~�?h�Â�Ni�Mz�Xdy��6[���^j#F0X�����Xp�2��JШw���.� �������wwLs�T��|L�'�,x&LFjd�9��%k.mG���L��?�����C(G�@qөŸ��ã��nf�{��ߌ�r<��9t�Cp�Ym?}a����rJn:X���;��X��2ކ���E��H+k���fRǍy�pdk���f��Ͳ��z.�;;;�9m�bϷ[�*����vj�fBӁop����=y��㹜�7n�7q�a��c3�p�����n�U|���]�gz�ˊ"��'Q�����ʖ�u�	��[�����ʕ�ά�u���\�{�)��]�Iyv�0��#-��,��wW��ܴ����K(KY��~~4_���:�\Nj$�pol~'�!#N��sy&����)��,=���
����)#q�"*��Ƌ��q9���N� ��G��f$o�Д��,�����Ɗ���dI��|���=���\�pw�s�^�.60�-����ptʃ#.g��i���6��&Ñ��BJv�����|nT���a��網�m�Z9����8Յ���Օ�A�4,�HG������!��g����8��u?&ikJl\(u�ߎ�<Ӹ�S]1gA���(�Ԧ�:�:�g�����?22��r���!�)��4�$y��G=;���q�b�1�ӣ����SX�2��~�����xP�)��u�����i��oa@HW�G��J��6*�i}p'?�:����Aq�"�P���Ak����U��Is��,֬�q�̻z���#tތ'��oQ�!���sQii(V��Xù����K�<F�"�~���&;��Cj�Ë���F@�ARFzn��|�8�mN�Y�d��|���Q��]�'M���k�����������7,�2�@���l3r<��_so-�/�]��0/�4�	r(�w��"�{iai��[��"r�cz�����?���a�';��ߍ�'�m�.�>5w�ǂw���x1��{H�iɽ�bgn���*��>���	���a�9�G.'�`N��@��]u��a���9���L�=	�c_�k������[�XyD�ٻ���*X&&&���c�ӹ�-����H{���{��h���=X|G��Dt�:�~�4Z�8�5dae`F¸���p��%��F����ö�/�"����˦�v t:A���>ڌ���N,gdkhح���FU��Ҹ��!�&�'�I�������g]mu�z}GF��k+},��M�ӊ����S���ƋŞ�S���"���f4-�������c��E��ҋ0�T_I����+�78�A�\�ƓƗ��F���b�:bsL;щ�M|ks?L��4YL�5��Yp���N�M ��ر�>$�yY��$��]�_~��@"t���L�������Y�k�j�=�q{Ҕ�������
�� ��|�n�:�d,]>07n�+����5Rpi�u����`y��{��S�0���v��տ�i�YN_oed��Z|  ������G��C�Q���`(�vVg�� f?.�/r/?��&�*�{Q�Q���N��5L�B���.���X,�XOq=][S3$�=O�H4�����&fN_�"��T�I��>0�'����C%�I�5�?ϗQ@��#�2���X�����VK, ���s:N�:em�[P��V��4���}���p�m�E�i,�"y�&9
X���Fdα(#TN�2��{_�vT�O�W0���D�?�!�)�� ���$�'�#�vd��4�:v�����qXN&M0���}n�*�_��B*+�P4�:u,9Z���-f�I�5�H.��(��$R�i�L��]�55+�e2���ʧǢL*���.cdkV.KlZ?����ـ����"I��r��!|Ov�㕦,FEw�XiZq���nޕ�i8^��uf�X揲���M�|Y��_kk�X�ce����I�zJ�wL���pA�}��3��%_|:6!h�O��#�&\<ރz�OZT��	��~��E�*�]0���0���=�J:<"���#�����M�*�'I�8,�i3�	/�����#�SW���$9����u@�h�b����}puk����hW�����i�������"��D���T���-��aG��}S��Q��d�i8�s/J1��F/�J����BN~�G��"D�E��R���7�5���y�1�;�r��u������23r�r�-�ɖ���O�0��ڏX{��Yp���#}��ǎ�Hr�&?��6�mF����J,��+�3����zD�.����8��`'z:V��K��
p��m�{4PLcEC��S��o �ѿ�0�
#��L� M�����k>��h��(��5bNq�`��?�P4��F^^}ػ���]c�྿��J�J�E���̣,����7o0L\ņ�ܴdH��0^jL�v�������Жg�aj5M�]v!�H��FR����}r����АƊf��u��ܿ���΂�a��yH+��'�r/66�	�B�=�~4t��8�(�ʕ���3� ���S�(7^���0J���@�%PomcD��{E�wj�t��GDV�E�=L���t"6c%ʾB�j'�<7ϩ1���\!�s{�;Tr�`�y;�n�u-4#���x �N%"�FS��d1F�v�GH����܎�s/n�q���e�����pҫ�&�L�M�E��")8�aSv��B��=�"���e�R��<��!L���
����|.'�`���c>d�򗋨��u=c3�����C�����Q�EiP���ɮz<1���r@0g|�TS��u���#��B����-��<�>D�a	�Jz��g2�.���{*-���8��*Pc$6�^�D��K\j���7�r9�V��hZ��B\����n�!%��)u�%�<��a~j8r˖-��ƺ{7u�#��?���f���閬�ŏ�_$�ӷ!�W��nU�dg��|�6�9\��4;;K��籮��]������S�å�8sN$�\����-���7H��=Oݢ��#�n�}˳�.��S[��KR��ʃ�H�}�F��-���E�����`���ݗ��}�Thh���^&�T�Rccjn�:����;�%�"�Nއ�zP`�I�J��ԓ�d<n��E���J�Low�n��?�V!�<�����p�SM1#�T�R�߇��QFM������<���/�c;�ѶA����%�7,x��v���k*0��m
R�4��#�aV�AYg����þ�<��qg7�����N�F�����ᰧZ����	�|�67[� Ȗ��J���\l�N\���I۝I^��@�;]��#*���(HY�1~�i��ao[��)�1�������mgtg]<<<��������9P�>zr����q�%$�wž�إV۩�j#H�-Ej�����h��᭑ɍ��h����0�ʶ����nwL�4����a��g���:~՝M��3�*�P){?��?�S�� �_%���+-u�]�oZ�z�:Y�2�D׏НG,xz��;���˺$����	s���[wy {Yl{�c�#G��]%���"�R����O�3� �)���*��Z,�WVGj0����9�r:�f�{!noo?����	(6l5��?�^UZ��L�-%T�v�bא�a���@͝��F�<��β���`�lg���:��3d��''+�#D��!G�����b���&�<��,��n���A�y�b+�SI�]�]�6���g�z��RW�w�� �D=���g�����E�	�Z�f�(�G�����ז�2>[�Q��-r���q�|�)��2� ˢ/>�B~`���S3��������H}>�P�:l��ۃ��s����M�r��{�8�N�_uU����ʿc����Ypb2��+��h`3��GGGw�.̌]�o��Cg���GO�Ӊ[�P&���[��TH(�zl�&�18�ǥ\H�,ҕ�w��&α��O��� b��2��C��1���$���M��3����;�O�ʂ��'�2B[�Jקq�'8��u�֎̎�Mr�/ہ8w���/�_'±Hl��Sp=�c{?1q9�X�����w��hJn��|(�F~�SCf.�ONVWW����"�xw�,���7�a0^B��_|���~|m@��H��_�(�l?lbw}���T�����!��`J\bb�)_R�ӱzU��~���.RL����;��'�[v��x���M+򖜎�"UCH�б����Wr8G�#��3�����X��e�Q��#�ӄ�P�����|��z���9R_[[��Yo���GU+��?Ć���-)�c|��1���e�@�*�c�\�֋}�_����gF~����]�s%}����� �䁿������
&6�����Aܲ��}�-r�/߻��#P��
�𰹣cz���u�/0��L
�א*�FW3��lUZW�
;�@�E�c��pY��e���6�**���|�I���ɶF��w��=#-��1�쀦�r,IC���-�v��Ӡ��q掓�YX��8p��˲�x�i�z�r�d�՝�";�AT_�	��*}ݕl���o�A�_YYi�U�>j0�D:ħ �Iw��W�`+33���?��oz��ca{�����D)Mߞ���>i�ل�v�W��X��"�3���� ��xEZz�8�P����Q��D�l�\7(НL���x�8C�5b���Q}#Kl�Il���d�]#P�ω�+��*�(�g�rn��{"�x���Gl�q������qq��y�%�ԍ���/���Tp.u�e0kF����k ��Z���E�.;�GX/x��0[3lD'�NJmȰ.R����+5��M��bܿ����}L,�)���cޤ�GS?�u?����������q1̨�1�(]RXC&��������/"�..�8�"g�G
�
Z��_�[~�[�1 ^�3j8^KR�w����Pi��[����3��:��=�$ �7?i�(z��J��!/��������X�����u�Q��tL�<0�Kb�M�`Y�8�e-�h�3��Y�`Ge�Hȋ�|k��ԗ�|�+�E�V���x1��B���]
Z)��'g'>��l�>�ý�f�+����@�g�a�f�T�r>8�w����Ϊ������b:M�8��ܲB�@.��?
]ZrsH0G�nf�����	��h�[����H��r��0��b��� �����Vb�qn(�@p0�;t���]]�ǋ�D�x�[��1l8^��u�%�8қU��ss9���v�غ�P
�0v�C�%;a''��N�Q��X����v9_Gz�&A�������N�@dz�y����m����g"E����
�O�>N}�.�{CTo�[�`Dgy�KǢ��^���3Rw�<y�
]0�e�䛪�-[��+So|�%�^�Z�҂a�~s�$�E�a��S�l�'[�����_��Em~��0s�{������xq6z�U~A������|��z*"���=�Y����\�;P��}0��9�\���O���˴�mv|�~t� �����>E�8IFU���*!ѥlq
��Ի���)�ФC�<���\�s�V*���1Jۄ��
:؎�9{�X�������0CV�/@H�K�4Mf�hY>g�����p$#]_�����),��w(�T��~~~��}���v�9�D.1�rrr����3�dIe�#���Ƞ꜋�U�\��Z��:���+��������S���x~��6�n�;��t���C�V�@�6��n�,��P�����59N�獀��<'����?u��~��� ����^9�5A�4.@ɔۆ�N;@\J����E�^��/���X�y-V,�˾����i[+��A��J���>a��3A�w�T5��ܽ����Ś�xe%ta�PT��**��1�؂]R���4�*�^��[������=E ��0�L��hXҘl�|Y��Vn0�:�:��,߉�����O<�>�s}�K���# v���.� _2�0������Y���b���\N��ٶ���[R�8�	,~3���w���ӧ	]y����+,�����\*���{�_[!���	V�A�D#�t�R0V��:V$��ô5K��\)�э�j�zW�n�u`�"�.�����F�9;���k�!��<5(�N#hA���a�]zN���.�����h��R&$(?!��%P�%蹲ER�����e��<ÝOW��$������OԝC��e�]��赐Wa�掋*Bm�;��^}]}�r ]�E.����a�dO����J�F��d�m�z�f �IL*<����Iw�V>$�|Ma�f�y��$x�����
�x�?��8.V������O�⥚{ʙ�J?+��rRAHxUG��T`.��8���@���2�]��'������G,l����8����2zFA��!6$vI2◴�˚��%�V�߅�#���ђ�����ސ͖�+6��/�'K�ڮ��]�=��6����_��~�֎�w~����^�:i�u�t�r�us3�d�οx	�kN����i�V���87$=��2���4?M;�#w��a晩8i���V��k{�B�$�V |G�B/&�Cݝ֊ۂ׼[ď���<���;5E��1��F�#X�V�p��x�n��� �U0"�G1�IUbi�f�;B�*j��G��4�'1l8y�G���'3��ݻw��<�K�/���Rݲ@_�ƪ�)1=��>ܕ�~�՝f��R�ؒa�|f/�T�n�����{�嘌�p�O�M��]:������ˍh�|t@��e��]^��V\�JX�Ekjj4�a�?@���VC$8�I����x�o\.����D�^F3��6~����T����g����*�Ż�����;[��?��b=�;H��$�R�:�}�9|BK��d:��]>������_��E�~��O}r6��k���<����IpIu������%f��\	��oPƜ=abbAӤ����O}2U4��yz UT�Pmbb"T���v�4�o�pg��N���躋S
�/�����ܼ�PZ��JU�|�r�Nm[��,�]��PWVi�OgL&_�|�Q
�����������H�}b�uf%`�\61��0ҍ�^a"WFig���[g�!��(�~(�d��&�š<'��������qa2J��g:�m9ض�^���`�-Z� nf'D�c{ �m�:4k���K���?�2[��{a���bǝm%�3�'�n<����w6v#H��SR���# ��7$��l�-,
�Di�e�+�(��O�U8qV�F��t�N�?߮������IB��Mw����n1�e���;O7 �7��c!:c�5@�1�j;,�WdU���������l�ա�O/X��<����_jQ�&ܼ���]�5o�ΡU-�p��Ga�t�_����Om8mk����?:l�Z�2��=]6�^@o�^@�>}�W�9	�����Xא7�'~?iVK++W���\eR3x�P��ZM��_��鎎��:�2�|q�Lr/���1߅�ڻp�)eca.V��Ю�i�r&lK����%�V��hn^���7hƣ}3"���槆Ym �����M��Y�9��i��#V�(~;XgL�ac��z��ȏ��9%�A�D�PQIccaf��6��0H`B�q� ����Ʀc'Ow����>p���I+��K2�ESOf$��.;,�iI�U�X���i�T�w��f�"�v��Hn��|�h�t��q��[(+�a�ڙ�b��W���}�&�T���@�������������C+ ���F���3� �B��g��\��l4�i�M��f���=��Xd��7��GpV���y��+�>�iy�9~�Ԟ��j�A����f�_))�o�u���!���Pjd�l��~U�Y��"jH�9Z��_ �8��<�v�!���\ΠV"	�İ�M4�]�M��BY�S:��0� $g�6�j�u�V+ss_'����y#���!p��܏�L321���rd�{�@ �=[AS�pp�A���ґ�MIqފ�F #�tJ��`ك��a�R*E����u�Te�G��Ə1��z�h4(�jy���g��g;qT�԰9�Qgce�0�[D�(bg#�G�T3��С=�Nܣ}��TC_a�`lC����u���@u�WP�b��3:��ED�_7��h��f �m�cP�R4�BZ�� �:^�8�1ɾ����~��9t-����S⇮Δ YK��VH'���wyGrZx{UNM�b�+�B8fL��;2?-�	J'�LT��Ha
C��Z�Z��d��� '@5w2�6�yTD%2�?70�\�f1JYY9�O��C1��4�wQ�lG�H2�n��4��zD2c�(��&�%E�XVie����h3%�����D��_�A��0�!T����C%���bK�AE�yA�f���MK޳w�0���	�D�s�4𾱮�H��
�6�%to419�5_l�u����6߿'tw"���3�[������0��$4y�U??{���|���p�@�[r��]��f�|��ڋ(��o]�u_����op��Ц����O5.x!�sP���wJ��N��L�cqfm2�=��=�6��Qs�1��03��_	��=�;��7�RH$�<��a�Z���ha��%����x~\��I����<`�;�����.Z�P�������oA���f�ji�A9�0�(��������S�>�a#�_l;�bp�����y̷ 5�ɩ/�d����P�����	;5�::߹�dnj���2��[���Vy��m�)A��Z=��/Al"�v�����MIy�����6�K��T
b,s�_w�ƙ��NV��B1C1�p��y����8q<K��8������y{߾�!H3�bC�c�Q�$��Oh��zz��Њ�|+^|(�h�M.i0?��
	��'�9�E�<���C�^D.vJ���Y��0nP$��D�g׻1#z�����f'��=���6��޽{�;_Rem��K�#�EE999�'�Kv =O�����#?]5�$�I�3���}�Z��-x�|�>��ٌ�f�Bu�f����˚��K6��&<L\�8���Ї>��nX�E����4-�>�~
������O��b��7~|�;UT�%0Cߟ$��x7wA%Ǹ���?���6��ט��H)�,-���]�o��w�PMA��4��\I�	G�y����t�R	� H2�)��� L &��.���u�q/�-YPu�0�@�t�K�����8?���-�PuQ@�J���mQ�n��`�b�Gq�*+Amy@&� T����c�X���ž\cݲ�q+��|AwPtn1��p_��&��,��Ү�
2���=��].46�g����Dϗ?�Z�)F��斖����>3�f#�+�dq���jR;gS�d���C�˺L��!&��M��Aϣ�-��P�˚ 1�&�-�G�+R��#��x�A
��@�	���/qJ$�4p��4��t���X/�@` �"�P>1ߟ�V�M��)D��g"̰z@򎘝o*§ �Ow�2�.����
bs����G���E]��Nl#p2���ҩw���i:}�|i�����Mz<5�D3�D�f�5����֞^�ꆗx�WT��P��N�������y�n�o�Gנd�[f�t��$T�Lw����ù6�A?l��R�*��*	�P�ܺ�?2k�K���m�JM]�RUi��}T	=l(Ů�p��EU�RyB��Jq���C��9^��8��l��&&���)����0r�hN�<������6}��P�7�����<�\w� �0�.B��`���cN��<i��Y�9z���_����n�g .��(#�8i��@��b`bSQV�hZ�����/���gB゙!��6J��'[�����%c��V_���� ��G^��PV� Y�L�a�0*�oo�8(
���K+����ʝY����\��G+��{-��[����>�_8�yY���Y�*b�:��N#;pT+,�ϲ�\+Г�D�w�s����aF<3b
J�aLUq�@7Z����r��T���L]��4*���@�7^֚,'�F�yGA�P�#�
{�bw�������4���O������1o88�&丮�&A[���������e9�E)����T�
����?�r�vg���X���c��82���>QCbs}�R�tf�F�����C6[�Cۋ!쬥yT�H��߅��z7�`cf6�E�=�����I�i�\�`=�9�>�0� �!�� e�O�ʺ-)N\wU	�3-�=��i�~G�����wԻ��Hw����|�X\�M믇��- �5{�x@�hF��"K2�A���|���\o�WA�!=m�G�u0&�v�>u�y�i�!k�60����m��,CH2N�]V�L�v�@�3�i��z��!��Zd��;���E���֡{�W��-�NܩZ�Sya�h��1=�V��EKu�glҼJ뱠hq2W2��Ӧ&����W<D�+�ɫ���/�_­��%B�'����I�'AQ�n?KI�����ܧ�ín��i��j�ÿ@�!��T��?dNY��r�
�g*GEE��B���PRe��ސ��؎�
3�OU��Bg�ʍQ�+�X�`�*c���VLM��}8Ӵ�� �z��mЇJ�03.?r�j�ҾL�8ٚ��Ǿ�ZQA���3�9&&в�� ����%O�|�_I���i"��v>w��a�έ��Z+��ǉr
4�k�,�ا�����|�����I�����N���בMA�ѮI))�'N(1=���0���l�x@T�\	���~2�1�Q���;{����jq��$��\�HJJ��V��pǅԈ��4���:n���$St� ��$�^��q��K���d��`R���i��{���,�� FP��V
b���k�fl��*AqU�G�:՗c���*�q��倿�"���e#�(3$y4���?N��U�6����%�P�������d7��O��)�����)$� ���Rj��q-A*qW���ʖ���&���2����?JQ;K����n\�n�|.~F��5H3��x�j�a�y�L 7?^�[(�;�T��lZ}���	��AO���st��J>EpJ��I���@�2�	�w}��w���[�C��/"��ʗ������t�ɕ�f���H�'=���d�N������/��kOw��%rRRFD�:��B�\��K��h��zʺbΘL�h>�Ŧ_�=QR���#������@�2�ß�N�}�Lw�H��%���hЛb��P�=ᙷ�u叐Aȋ#����;��))~�Z�GosW��ĺ̝���	r���y����Dy�?�+��⬜�� נ�%��̾_�✍̣�!p#O�^�� �I�h=�%vwӥ�X���G�� �� �EML�ʰ�\����IJ
̛��%�5s��t���uQ4�i'��Ȟ$ٙ�����0֙��	�k��FyP��L>���h�_(j1�l���=�9���祑�V�5�<�>}
,B}�^�Z���u�K8ͶFh\�OF����U/�?��%�0������z�T������_P#�P#b{�F���n�:�,�|̄�KҾE�GJ��ZU�yȭ۴y� xL�9��.v��X�Ƈ��wϞO��M��ԅpi����*+k8P���q���j43-��;����� g��c7�[�`��aE&��]�mztz>$6i�b��L#�����Z�~}d��G����Ld�?ۄ'&݆����2��7�`�����F�c.~��:�>����TVv�x�����L��E0���U�q�U�8��*A�p(ά�b��"�hf���BSS$H�����,	
&��7�r����^��Vf����!�}u@��w�4��nˁ��c��u�SRZt�{�<��]�M�tm���!HS��a�'����>!��=%x�~�p�^3�=�@�U4U��u�h�wz�68�dvD���
:r�-�}� ��M��\������*2�Ȅ����*ϩs������璸Wg̣�ՙ�l=(��l�+bne����A�KI����n[��qJ�d <��T []���5��!FC���NW�SG�Z`���VP���L��j߽��E-�=��F�ԩ������;	��,ͦ�_�j�wpp�E�������y�<�l��Q���n�D���Q|�á���G�2�����U���������L)ȋaDD��b砍��T!�		yS<�y9�h���~��H��~��]��Z�B���k���������PQ�L<��ј�tO@8Y�����*m-9Ş��lZ+���y�!2�gW���-��W�rjbe�[e��~V�7������v&w�z�����u�5={�c^3z�p������SȤ�i��Wc��@�0�E�ľt�����@�/@'�4�?rT�T�����M��ږ��w,�X�QAX�/*̰}�7��7���*�����4G[D�AЅScZJJ����W�(�E>Q�7X���X#[pټ�͎Re�k'�wz0�R�����GẄ́��xeaL�4ڌ����o��S�E��ߵ�f4l�Y�a���K$ɷ�܄)���W���t�ڶٻ
�y.�VljCdP���^:��z��������Y���-<rE�$����]�*!�G�/.��L�@ؓ�ϚH{�����[��ų�E��-E)��}(���혪���ﬥ�K��&����2΁�h�x�g��������叄���xJ`�V��~(�C�51�*�k�wZ����?��49Ȣ�v�0C�3o��F&S`����p����|_����P"YU�<M�y��)W��d+�!PTT4X�U&�8�`F��"lq��YN���t'���+ٗ0���4��r�k#�&ݿ���~��)�%F�����f�����2ݽ��_�!l��2zKZ5(>L\�t'A*Fy3iy�Ϣv�o�_W�&L%�Q�SS>��	�Ջ�;�<44T���ޡ?nbRJ��mN�G����"�/Й�0�;q'd
�3p�?X�5)�}ъ f�n���n0��?�8��`��i|ѭ2�U�i)�&CWQu�����p�
�IT q�������ZN(�q�u�P��~(ï�B�%
��L�	#� ��OC��|���J�',$���w��,�p!?�V9���v�-B��d�3&^g���<P:e�;m=F2&�~���3)+�Le��A�liav�{����	4ii���hZ�2Vx�S�c{��ܢ�E���Z���+D,���ՠ����dr�n��C��Sɱ���h�[9��h�M&+��~=���X*N�1i��)_�Z@[z����/q�Q�h���2�[%)r�c��'�X�����A�� �3x��`H=�U�
c��/�����DJ��߈�?w�}9�����.���M�w��H���8m��r1�T%8��)Ƈ52=�s�1@	pwa���K����#���+m9-�������F�Ӷ���E��Ϫ�a+��(�R8f011!�9d�F�V�re�0��+��3q���ae��yn���k�Ѯnr;���M��nǝ�*;�������U�K״X���lM��f�=i��m���Y�x�V�3�zO�驞[[��~��l���/��y��Ϗ�,��O,�\z?�·�X���Z�6߁��:p��������D՘�ªtč[il��ol���~�ܟ缼r�W��Z�D�V����2 H����a���(M��fd!�@Е7�����mZ���0{-���I���P��k!��/k�MfTB��wB"Í��8FUEق������sʉ�5��Bp�֋����7�d2�#�(��#o{�+oo�9�q;�+����(�0u�f�-��q��{��)���}�S�5Vs�3>>>/�������y�ɪ���m�/� u:O� �B�SRX'�s[�x���MK��ah3NU��٘���<�D�*�
{�h,������C\4v������ـ:�5֚c�F���Nb�����T��SZ�.!~��8�x�>���*��ft���E��+�}OV=��ý�J��b�.z�Æt�pP�|_�j�7�*�,��=��3��_o�N�ѝ=9�?��7{-&����S:|���T7)@���J:������N�i&c���7�pDW�������,���!A}Q�{�(j/��$�py{ ��k�E--�լ�j-y�������?�P��R�����E���xˣ7���3 �z�ߵ�}��ֶ�H��&����Z�����b~�f��3L�z���_���I��v`���ev@�?���Z��ޢ��F�~$�ή����s9@[�/����%A�Ci��Bt�|�bY���|b_շ��k�G�B�rQH���zS(����p��@�ǅF�*���`�x-d�"���ׇ�Ќڱp���`]ʁ�Z[y�U�0jJ7���59̌+Q��2�R�u=��u��_�+����֣��t�,d��D�|�_��b������Ǣ����%���K�����J�9�)$�q�>�_�oE�
f�����\�n�ղ1���ӓ�²�(���q�&&*Z��/����0y���B;�s� ��6B���A���c*���L���~�l�q�G\��f��q��������/���Oaw{.I�	��,�'g/LF�5=������8�q�a��+\�I��Zk�;�s��]���-���P\"��Qo�w���~4������틵�O�*��lh@(P�z��6��#ե��Ԕ�տ�I�D5�ӥ~�z5l�#�PY��j�O��wT~x(�G2�ɫ����}4��U��_^�bd5Qzٖ�U?�����A�-'��UlI�g�vO2�{����������0_q|��{���-�㣱��#'p����ɔk�~��`��jq��掎����#8���d|�B��w௛[EE;���V�i�d�e��-D �M_�B��G����_�����7'����GB�v�vrr�O���.Y�>�Q.���p��f~�ZVQ�{v������ċ!8�2��Nz���?'� �QU}ff�-�}{�' ZM�A���73/hfUw�Y찆Y�I�60R�&���(%���Z�XP7x��������o./\���,����a��B�u�Ӡ:�U�bly����0�����,�О�k��?%�` �o�6�P����g�0��r����a0⏡3C�I����I�t�z�������{o�M<���TT�>��+/���0�)Q(d����_�En}���8Ѷ�[e�?�����Sأ�%����0+K���|J�F'�Z YJ�P�9�))�������Cӓ���k��s��b�"�M��Ԓ�_��1�&�� U�H5{�
����#!o��U}�Kh+���R[M@��H���*n��X�q5�'���#Խ>4uB_P�G4Ss����9�u���N�N-Q�ج�Nu@��é�&Z�V�T5��P��+qCb� =S[�O{j����"���g�>D?J	�M��K->ר*�Э%�58���a@n9I��$K ����������\���]} ��L�g �p��,���&RQ��g%%�Ra�ҷhΫ�=���w���$t+�c_�d�5��ؔ�A����w$װ?)CIŁ��Z�K�+�m�PƗ<���_B{�07����#���7�?zN��f�i��Ȕ� %BF��1ȄE������_����a*��I�r
�|�Σ7�� [%(�aά`�T�*h��g�i�u�z@�R���JZ��W�e]�X~s�8N_���IDu����.���pJ?����ց�ǐ/�QpR��R���TU��<�Њ��G�%q�`yK����ϖ4�JAG�2��c�2���l�Ԕ�����ZW/�z���$�u ��2B`A]�G���?��wQ{fU8��mڵL-��?��ي�_@�"N��"�8;;{\���-�S�)��{-��5��y?� M)U����V����T��˨A��!d�i^��Pl�6��U��a���u���p���fe}̣�g����A��(w v$Ju�V��gV����A����>��ְE��>i<wU!�<5e�~�
����_M�):���AT��4>���Q4���8v�$W?F{9$�����s^K㪒X�":�x2a�S+�&����Ƥ9�y�Z
�0�{����*�Z��A�bW�0
��+y���[�t����7�:�!֘ś���O� "��e�1<�dT����J�s�KH�h�[EJ�V�����9 q�����b5ͬ^I*��t#(��Mmk�=m�ZUT����}C���� ��i��⎆�BW��.���ii�@n _D�:�)).4�՜Q��KJJ��η��(B� (�ܙ�_ ��e���M�H����/�ُ�#Y���|e�֧Ub��0�xb��dǎ{��V|�P*#�u��/�o.�TJ� �q^Cj�Jk�j��G5X-<�D`�7�`1kQ���.��z�ԺES_�Z���l���|I��(d��Vq�� t� ?	I �KVUk��[�5�j
#����w�#��������v��0�}u�s�W�EE@a� �s�2��ϲ��U/��@<CoU(=��İU�w�fb�	�(�-�q�Iˤ�v�/��IP�������^/�
%������ͺ��d��yn��Ⲣ���_@)?��[���X�]o�d�,W	�뻅�����H~O�� ��ټ�K�w�Q����:�:���Š�������&o��s�Ϲ�B'�I��Y�N�B.�TWU+��A��˹�7iޫM���1�bU��.�*��P�Ƞ��Q�+��`d���wD��u{X�6//�@�\�3_h��	���3k�Jͭ���BFW^񃧚a$��-�~Ammmŉr��w���D���W��&h��
���928U��wp�i��-���U ��w��5��QUN  ����|�aD�����V��{��?qf�Ui��ԯ?� A�����sI����g�:�{oV�����
q8�qR�Q"E�ѱ���th�T�4���&�aK4��ٕ� �L#'M��JE4����������{]����k_��:g=k=���_�}���+'�(b6�|���O�>2 ��܎��$���1��ʪ{�g�= &�CE�yB��'�a0hD1@1pܶ(6m�����L�� �0���h�/?�P�5�����K�,�f0�<���Ŵ��)����|�\P ��C�lon}K;�������1;�lY1�����>@K�#�M���#{����[+��#ߗXURQ�9��P�z�t�mU^����]$�'�YaPE̩�[jY�ux5�3��T��KP�5��׾󖑒G�KBɭ6��y��G��^����"�3�++�y ��0T1Ӧ�TB�u�wi��g����0��}�.%��`������� /=z�#�����=�v
�"�;�~9/�����(�D�Uw��)�T�ca���3B�I{+���e&��^��a�1����:qT�4��عs�2��D1�n�{h��(�Լ�����`�W&Cx&�CKQO�MU^"�zr�G����`4����˗�C|v���*���ދ~���}	=�����JH�ܺ�	�,<�m~#}���.��RrJ`ͬ<ɖ�4N���	�{���y��ȓ�3ؗ�:��?-�4���{�� ��cI<��fx�k+B��޻���O��F�]dXX�4�U݅#z��{ |��H'5� ��Qm�P)���c؜�t������W��_�tT�Ks(eon.��QN����}�W�.��><h�N�"� ��Ĭ��-��s��M[���@�* N=}���a^r����/�Mp-��k6�}?�:N��@��Ym��^ܴ������8����	bP�zx��1�wU}<wv��F;��CrT>g�n�҇�+���M��*f޻����Q�V3��)U�@CQ�`��ޠ��<�W7��x�.&��A���~�\�G�D����I-}� �zK�r�2%uV@_�QN
��������Yț�g9Y1�ƶ8
[�Y����ԋiD S��Vy���[t;v~�X��,��2Ej�{zv�p�,M50,kU��T���l�[\�3)@��_�H�v��q�������&��8{JQڰ{�_/�Z18���`�-h,�ߓ���9C��4e���G�(h�:5g�5��'4,��MI}���TgH��&A|V 7< 7th)6!��T�O]U5WIO��	8k������9����Si���,?{�st˛�I��
j��5F��������~TE}B�*�-��������F�O_@��RXcu���}�b(J��3�:�����=y��Uq��w�9�\�t,N%�]��N�f����T�f�1<U�&t��=>Ҹ��ջ�egM��:�u��T����5`�o�$dس����D�3fY��:�&0��a>X�L������ς�v8�'0	��W�Yn��wf�������],
�.�*/m��Y��h��s!��(8���F���#{�{��=�m3���O��7�bO_+�ڱ��&߀���/��W�F��51�o�����g�����%x�K�����/���bjyM������z菙��E�V�n��-�GZ�߬-݌~�p�]b�.D� ����n�ʻ��P3�t�����K�w�`�c, ��"� L��y�4N����~w���P���ϱ������b����߇`~��z��	�^6DSL�4׽�ҷ�����(���8�� ��X21\*�����`k)hF4�M4Lu����+��_��9jr� �Kw�n�J�I$
�xz?�H��]�t��I�(t^���Y�Ϙ�i�-�n���G�����79_oQ�o����e�В
�/ߺ�����?�+NA��&�#Tr,�O��Z�>�%��vȨ;�߽a9�x-�Z�e���V�C��F��H�V��-�'���ܖ����ؔR`Z%�����s�9�X��߬p��G΃\�g�߰h���`�=��E����G{D�##��u ��?�0�A���ܦѪ0X��\����%���	X�ϲ����zzz�k�~`�^�	��ca������Έ!���Qg��P�J���� (���08�{3��<f�^l�5��fØly�4Gm�JMG`.l�����*]�Cq�e�:�
Ϫ��"0{%W77.���!��gS���C����p�C��;t�>�$�o�j�TeH��Q����������~7�.��J�Ah��Z�>n^^�{gSb�B����uu�6�� �ԟ �@�wi�
�KN0���A@�B��1��L9���0ם k��cx��z�Xhh�q�ë�r
�H'E-�r��B�>���)��ǈD�&��eľIuG�V�ty��Xa�Sgbr�443�=�maO�Jc����6 q�G�4z�T�'-Z�z�2�=o\�u�leS�7�]%W���+����<ک��wPʲ%�ݓ�ij!o�)��X~#>TVA*g��c�P3ѼӶJ�K<T#kƌq���S)�����8�X�\���%T����Ӑ5�ʔf*U��X�� 6(�������4h�l�a���@�(p�ʻ��?��J���+��)�(����>[�uO�={�&)>�@�p<�>�Y�Nڄ�es��ra��k�y=b)�T����6N�C��I�y����#�~V�f@w�mZ��֖�x����яOT��{KL�ZEá>���@�1�3 qZ�Tʰ��W#�ӂ�A1�Z�Q�rr�;档7[^��D����j�
�F��)���222`�5�v~��'����=MBU74$ӛ>a��D<-�������t�2;iZ	�� Q_�n��&d��.�x���ߢ���L	�e W���V�pȷ9e�bp�.�Ź�n�Cb��z2�Umj8�P�&sI��%WgK�Te/R�_xڌ96퍂s��{�l�����\��J(�����s[��U��u�dA� �E��ʅLIoS��zu���1�okjjjk	;e@V�u�aG��#�������Z�1%�{�9�<��,:A��4U�@�{tX�~o��{�e��
��|j$�[/+�#w\O�i�\�C�k;�����+�t��~ݭ5��kw����@��vS�e~�V=��^�z�ǂDY�vJ��F��×F:~IZ-Z�gQZV��fJ�J���[E�N�z����b��kJ�����~[̾/�`5�q�7�z,HLjt"�'t6LO��m��$�]/;� .��
>g@��?m�*uX�|Z�D�������@N��[�QՕ�ȹ�/�pa\G��_��a�o�{����ׁ+�ˎ���H�.j R���їPVr�޶R�����	��	uGn���|��8�����<�%��k���>��S�	Ҽ��@�8�.���Q�э;���k�GB�T޽�А��u���gb',�������n4e��:ڛ��4��?�JZ+�}.44T;݇ؿ���bb�/O��Z�=��x|ݑ�,ORLU�G��tm�Uo�}��V�ז��^S�G���}�"��Si�ND���:�����a��S��:���F@�:�e뵙wL�077o������:�ݮ4mB��y_=�}�h)U��%	��4~���g�V��UY���W0l�T�����Dxk�����q���)
�w@azxA�5��C��~,g�G7��en�'�p�Όm?�������L��֫���r�����}�}��t��� �u��Ei�f��ɧn,�?��A�+���-H�q��sMwR��q�º^ i��d�B (��ը����ő��?�'Ц�2~�#����ӧO�J�Ę��C�����e'��� �[��a�� �]&��
xb�AP߫=�ȫR���!(����;wС���+� �U��В�h�E���S����d؛���<[��0��S)+5��2�������e��Wև#��2�#L�N�K�*y��D6Jz�y��
]�2��l����ë�����ɜ���y�����{6���4�"������ �C-�_߷����D�eM8���ޒO)�c�^o� ~ў5U�A������s2po4�<4_M]�k/6�kX�)��F�_?���������⢯��Ǳ�a]�{H+Un�BǃWT���5�|+���ePpN�J��'��v��!�Q�4*�lV2>pYs!lg|�b�Q�k1��:E��*�btz��q�����A��81��O�����3�E���YI� U��n���^��� ��VSN�p�>2�^�}�1�fs�����K��0M5g��H�.gM^S��|Tq������y��t�O>5��06�͸'��)T>�����W�F��V�'!�(�ׁ?q����$3�M�7޹³��j����|;��{ 6!�9��T�gJ��h�4i5_�1~8c��/�1/�]�,��!o=&��=�ϑ���z����jd)adT�;x�Rpi�۷{�jI����3�3f����o�?Ĕ�D������[�#WCZ��v���&/�}��Р)(�lƗ�V:�t)k���a�obX���'/�^�&��f��῝T��WF�i��-pf���o�=��bRF�Q�o+@ҽ���Ӕq�9��+�
��%�������_hC3(b�tᆇ�#��ݻI!�	u�z��D�@C�m=�@=�d�/�gq�P	6�\"����O�����&���l�-����Oŏ%�gp,KӨ�g=\>	�������������<9h��8.*�A�&�34���Dv��JJ�}\p�\H(�
�2�(_A�@�W$Ւ��UeQ���`/��T��8����ax1��MhR/�M���d��!Wd_�|�r-P�
�li#��ͦ� ����%���+�rG�z���R��eÔ4us�K��U��m�}x���jvs�i�"����
l�Q|��ZU X�(-P�*����&���$pX۝J9���������������;	ԭ��.��lXX�6��ʉu,E�h_찵�y��z}�	��d:4�����G���A��!4�̫6f|Hg%C4�^Y$�z-G!DN��c����t9?c���yc}|�L����/��lA� � �ڷ�U�~mˆgr�7���=�.��я#/�����\}l�� Ȇ�4�Ч��m����ZE:��k�7k����sȶ)uN،���8o��K�,��W�~3��z�"Aj�y��8�)��U��N�����W�����O�U�W^�U��;V�G'C�����G¿�����?�щz�sXj5���R/����1��:H�����X����tm�o���˷�a�#3�S�W�����r��qSir��+V��{�X=���{w��|�+2�\�����P��c�M�C
����:hq�`�碯b.:W!^���8�O� %f�"�p �.�����$&��{������D�W�ml�Zd����֓�cg��f�������~^}�|����_�2Y�<Z��ƮO�����WQ���ͱt��Q���� ;���M�g��y]�;۱� Q;�]=�/P�8x����Y�vƀ*�.�ˀI:Ua��̦b@;�fk?�����V���Y�$���Pg��At����.q]�-�-
�	v+y��(O�����
8���JRz�.�Q�qh-"����EEM�d�I�`gC�ӡof����1RZο��D�NUG�{���Q�9�c��Jo*���!Ƙz��!S=F����ULaTi�]̸�Hn�}�*�?���dy�u�?��G豏{W���t�ܭ��~��&M�ry��P�������b��l�
��|�N�D�>/P���%G���j����4��h��aGΦ��=ik��/��#����b���p�C����}5��'Z�PWGB6��Pd��	[/�U�<�[�Ro*b���N��`Y$�eS��$�������v�&�ź���E�8�(Jj?Rv�(̭��R)#R%��C w�z�Q�c:�G^ڴ��4���`A����h���T�)�ވ�w�K3e��Ts*A�N�E���'���p�K�8�����l��8w���w,pC�q>v �֜)Y��E�H-L\���+RO��؏�.'���#���cXVS�c��0��w�v�+�!����eg(P^� Z�I��,h^I6qD�<x��H��@���·���� ��n���;M�U��>9#�@�oZV�`���Aϟ���G��qF&ٱ���v�]JI����Õ,�򶟇���Q#z<<�k��RT��k�؉˾�e�F�L�Ìv��4QD��A�\C��g��1�te Lۄ��__��X�������\Q8K�{G�?��t0:M���k ���s1}V�Ӡ��0}*�-� ���XЬP$踤c֮��0A=�Z�$4��p�a9��j0Iq*s'�*�6�#�Sn�j {6���a�n�`����Rc!��������.c�h�F7c8���Qi�b������L)Wu�N�<�>�T�E�&�YA���06�@�	�H�U&M�OOs&�`��3*�ѕ^@��E�4��<\��D6�':�Klz�FL��P>OA�>	+�=�+F�$���p*��%��q l;&,v�	X��LrB�/�S����I�`��`c4�!M�x�C������}�tKL�2�ś�����"O�K 7�e�,��#*�=g�Q>�Ng/���IH"4c�߽�N�����TAZ���$Ӑ��!���UNW~{�
/j��t3`�q���6i�`j�D:Mx_Vtr�t�Bʌ/�~%%����E�qR!*���D�����XD>V&TO��=2���#����-�
��>�x�xL5PK2�W--�%�(�w3��}����~���,%��4@�Bh<ɑ��*�63jleAO����D�q3^Y�;�K��P������;_�W����AM�>���(,x��X4t]���	�]�GQ�ӝdWA1�F��xC�`ޜ�X�k ���_�,��jH��@@��b��w'��S�*��;#��;拓��,x��X��z����ͯ�yw0�:�����ɔ�ג�d��Q}7Z�۞���W�)X�ryĿ�k�5w��VN��-��>�� �.�B��7&�7'{�;e�>��ZA>�A�e��U�{��3� ��N<������D����=�B��L��.n���ʔt�Leq�W��Y��-s�X���K%0���B�~y[��}�=���={Ǹߧ*��;D���8��:�!3s!��a�~d�����μ���3���4a��V%gS��W}"�Xz��3Ċ��SicxY�7?���b���!�قXs��H:��}���}��<�>�7^�emN�A��Q=�Z�m��
��Q��=sӖ����@�Zx�q�	Q����.��<�������/-RD*�݋~��_#���7���b7�t�
����;|w�
Sr��٥k9�}�!��fB)�Z��p�u࢏�{�'25�p>��Lh��A�E1���s�\q���1�ӳWeP�d@n7�4iźE��h�U6bn<����� �C�_N�84'�E��;� �OL�t@����g�9��VnD�g����1����t�C^�^��?��OuO� ��ga*(	�8����v�i�Û�
��Uu��K�s�����MI�����^�M��+���R�,dNīWS�������P��8�58p�O���l����L"����K~�V�z%�VT�ρ�U���F�_E�Z�.쉈��|$��1٥k=���,��Pr6ot8�fR�\br�ө���c�C .�7^��Ÿ�cN>����J<��?��.�It��f4�'f� 7�8�$5�86��;n@��fmpQ��{=_�������n�(��*h�టő؊���?�w�J�1S���D%�4nޓL7�*��mY	Bg�S���$��=���{nj��?ò�"q
5	w@l�Q��-[�*T�DLcH�v������I���	�h�fg��`�>Y6����ۨ�x���c�81�?��u�(�T�����}Ζ��՚�Ȇ3�πJ���=K!
��?�b�l?x���ճ�*��I[�xӨ4��e�A��*'׳�)�x]h;I�Ɵ�g�vy���+O��N��VW$��i؄�y����=��> 0u�J���.��A�z�EXlq��Ԁ�bb̵�i�bl+����r�!�U����O�8U:�w��OÁ*d������� ��+F�G�?�D�s�
͊Z�z�dK��ȡ|"�����*4ɧ�V|P*`����3*���Ah �����Aj�F[��(� 0�zfAU��m�DU}s�S����B�����|G�{;7و���E��g)RUMH,m6�oH|2+� r�������A�[ݒ�4*�1���Y��'�zE�c�ޡ2���6u�QٚL7a�Gn�$<������~��ДMG�?�^���5|��<*�u��� s*��!��R�@�W���
��? �y(h��9��":N��4S�R�"�|�y�5�����v�6�y�]�� 	'�gT�-k�%�H�Z�M;���TBK��݆+����~��p�dC�L�x�yd����u���F5s�p y��N�v`[�R|u�^r*�����
�
5Z�#��:v���7�p����D��� �<�?�Ia���V�6�@��+&��`�pc�ƴM.]2S5!S���ֲ�Re��I<9~P��"��1�R�w�J�	L&�v�z�0�r�ߣ��3���9�m�8�I{CAl ��t5��v�����D�	�:D!�ճ�?��w��0�q�EG{U�6kO`N�Qw|X0�c8g	忭�Q�܆)���>����G����g��\�N�Oۃh���s|�@�]�y#¤�1��?⭌c5i��^%�y��w��ã�'�=�{��s�\��̈́�ß���A�\��B_���#Br�`��|�a"s�U^����`�9�ZB�B�S�H!���}j
t*��Js���S �.gEW��"�
��n��h�����5&0�r3 ��U�Od�v�n7Ű�O�^^�+[Nқ�Z�*zݓ�ڏĠ[�6�*��H0�΅��]͸Y1M4��2�5�(B�S�<&�Ok�p-���У��Li,:Vi�I@x�	�c�5(:��xtS�D�Ux7�(��@4 PȨagVk��?��1�~��%��d�����TӉm�?�0�J���~���wa-�8K]�-�
���x����ܣI��}�TY�eI�](��<{"#'�l.uwK��I�@|�\�.af�-4��C�8T��>�IG*K��fI��CxK�j�n�Aj]�?&�6�b�f��4���>|����N�7��d5c���T�wnVP�.���0�r��I]gt�c!	�q�N�~LtL�l�����H/f�XbR��]�Ȕ�`���t|	#	ӛ�^��7Kt�/׭�P >�k���-�]7D�?�M��i�L�:�5
�kEi�h�1 ���/�x~���#7��z/����<�H�kD���^����Ɗ��q�lo�!O��lap`�"��i^��MB��3:ɶLj���LA�ʟ7=��t���eN�;Н^1�	 ����{oy�
�gB�ʶ1��.\j3tk���~�3Ҷ��6HtbW��i�넅�ؖ�D�ZnE��.�ע��#����^|LxD=t<5	Nw�)D�#�H�}K��Ge�p�� �9����o��푉��Z����u^,�p����� ۼ�W���D��Ut[X�
d��FQ|]����)`x�Z�]���W��v��&E��et�����Ҟ���e�tY��]�u��9HTz z�ʫO����Q���M�o�f���s(��'��&�
 �u�ɛ����+G<,MV�e`���c��iaw%c>{X,}��%ů	ܝ�'w�-D����q�,o|q ��u�X�'�x��n�sJ��>_
}�n;"��O��K���m�z�n������,Q�5��OH��:{{{a�����fO!�PWAC͚�ر-�҇L�?a>�C3L��VVRF$6~�&����T��M���-4""BhB�\C<4�����x�C��D�5�GX���	0?��b�`1"�Y�;x�XB慢T�QR�
"�	30^*aD�x���	�(�
����,A�z�P2��R�Tey�����:�ў�t3n��H��L������b:����²a������#���#��c3�Vm+�.�ygUƩ%D��MI1�k#����� !�("��|�)S,4ޫ�AN�v!�{�t#k��װֳ�8����3�U�nD.��kz��0�朧�/�m�T$Rz�,�&Ye`��bx �:aÏ��?!Yn;|�R�0��y��-)4�,t�y���P2;�`�GM�(@�|���t8CQpW�x�\yV4$��D�#�Lÿ3��]������I6�{ў��r���Y�<���Swk���)�r��Y�AWHę���G�otP����&�����/Trfi<Y //�?�E3�txE�Q�v�¦��d������fF�u��U]�������&�ֹp�cݡ����I�/xpp���=}j�u�ⶤQӢS ���1�`�$�p�6�Y�s���;λ*ԅY���3��s�#���6���\:�����@�!g6��D<��+k�w1梌J|6� e��6�l����U#}�J���'C��9ɝ��Od�b�[���p�'r,J"�'P��1�;b�UPc�l���5c�d�&sn
�r�էu��ߐ�3�V!��%X_۟`H��"�*p���|���U�4�ү_�l��u��og�y�&�S��q���,	�d�-��lr��}�@pˊ��z��Z�B}����=O��n�|ɑ�##��oE�D_��x6{��A�q��]�r�W�_A,"��y����D�Z$U�����2c:2c�eM{��&��*��VF�r��� w�t6_}S��eM�y�'��	7�L䏬L{Q�̇�n²��w.i��_�e�L�a�,���$
��`�����E�&!���߶�?s�o��ٴ����3�D��ӚT�6���q�/�$��NPFEؼ pg)���
78���K�����c0���(�Jߡ����T]ڧx0�ݪ"�W�j]MCW�(�-C�;ɮ5=�`l"��;lpg�ֈB���O�P��
	o5�gA+N\�y&�TZ/��yiฮ�E��@�b��0��*FᏧ�sf�LCL��S�8��&x��
Kǉ������e@��96jo��JK	V<3��f|��`ϭ��=�=�mB�>�������>�1G�o�M�Sl�$��Vļ׌
8*pT��Q��G�
8*pT��Q��G�
��&�A���!�?2u2v�[#�.@�9��a0����
�r[V�gնN"vۥT�Ƨk�����숬�I<�k��V	»I�U}<4�%���Ph4����3���a���'�3��:�1��m�Ɖ�*)��ya�n벣��cA���F�_9R>o��O:a��fN3���#8*pT��Q��G�
��M�u7����u�ʨ�8�tj��gi��5�C�'��bS�j�B��t�]�'#4�2��kF�
8*pT��Q���/�;VI��'N��;�r\���6pa(���}���/���{_���ˆ_&ұk�r����I϶Wyy�*��V����'-]�b��fuE�~�qT��Q��G�
8*�������N������3}K���u�Wy������d�E�:\�
�^�Ou�<���,h���sg�>��8>B���c|0*pT��Q���g
H��v[�i���Mgf�\�o��E���f��ݷ��_�:����ە���n%����Q��G��7�RHV�CA���z��Ik|v���9	sD�=���Ï�.�-�۵�Y�� r����"Uu������8*pT��Q��G�
�?A���M�c[����=ݓ������U�08�++��LL�4�t��قW tT�$}�A?�իT�+��2_��;�6B}���
�?O�Β'5��R�e���. x��}L���;O�v�-��M�Ӳ%T��J��}�j��+����Qp��D/�}"���\.�6����C�G�����/��9�C�\W%�ֵ{k'�Z�醽�O/�Fm�b�u|�k��ư�Z�w�������O�b���oj��n��b�^�e�����V�_R�8z�b��%��u�g�WQV>x6q�ܜ�y�Ү�t�m{�:.[���sP��iꍡ�v"sf$q�L�K��_����_���XzD���I�x��f��px�:1�m*�o�������q�=��^�ރ��t���W=��H䄺#�u��e�p]���	ư������Q�]�Rʤ�cE^�I�"�8�WK�O�6Qʛ��L�	����zA}w�'�DK�
LU��*v�����KG�e�I���hH�� P�}�׃_v_�H5`�Yв6.Gۘ\=󖄅���'oo������}�_��.6���)�a�G�,��k�+/�/)�����bob����2�V�N��Hsy����o�n�Ϫ��Z�Rw����M%2�	�^I<�u7���X��{�9#�Sy�f
Hx�m�!�0V��fW/c
�*�E2�WjN|�k8q�%R��
{�f��|�{;�vb�iq.�����_E�M؋u��t���8�|mX��՗k�b�n���5��pq��R?=�� D����n��"[<�ŷK���Nb%H�]���؛��-��jY����;��W��%�y�(}�U�?ћ\�I�Xsof�ߟ�7��H�n�Ih��
 ѭzx ��@HҲ��>�}@bí���s��^5�/�3S�R!%������jwn��Nޫ/�"<��9����9ɞkH��7q�^Xy�p.n�*��R91��k�~���B�/���"������M�77S��� ���|�h�0 �̛��zl��:D&����)���Hvy���Sq(ZI��2�QG���&~1���N�Ԑ���.��)���g��%̅�I�;O�%��x W�������i�Q��M���2�ݫ��i����
�o����jF	���r�����]��>oc��k��	� ��IuIj˕!c�� �XWy�˒�3nΌ���}�A��#�<�r�<�$�{��72��IY�����ͅ�m.ZIFo�_����:�ec�ӷY���Ϸ�v�~e��B�g{��Kwwl'W?���J!Q�&��a������ꄕYMqy�����]�m�у�Je���/��al�uGM��r!*��L5�K�5~�v�7�D�3ҁ:���/{~CI_���j@�i�z��6%�@�:333�MɧQ=Ʒ�\�eP
~W�w̟+:Λ{��j�����2�iݯ�������>���P:�ɡ�y����!3����4�++�S���{��+�J3%d��}��6�#e5�B鉄�f*r���_˗�������]]�j���_a��O�a��ʜ8������˜0��,�&�"���¸)(����ax�� �\ѯ�4�8R�J\��e�L�&s���rb��G��ΒXv���;�{�{ ���Ǎ����'d���:���6��7����!Ҥ� p_�//л�=d��s{��W�&;F:�������w�[�t�iY�>��y��<|֎L�+�-�O�/�������[�Pz���(�LE���D���~����Hʐ���_Z��R�H�#c̫�RLFPD���@t@F�_\�m;�j��.��䰾��aV��;���lr�\Sn����qx`��\��h��Rԁ/`��O][[[-R��oΣgb9�դ�j^��q�|�?®T�Иq(�u O�mr��,v���b��u���8DQ�g�;f�$Y�����G�u܌�.��9��79_B_��I����gӠ�E�j����ُ��OA�j�#��]�!���G�ܖ�]�T�9���~gPLs�={�{Ŧ�5�rv`)D@�ʛ�@jUdf4vb�<��̙r���+'%Ȳ��$K>���d�9�8[�=WF�H�'&����v�s91pj���\1U̫��$��h��������:k��O����_ �B:����p��dd�+ץ����_x���ЎTA[�w�p9s*�ر�h&=O�n~�Kn��S@�8�J���7�YY+��nr����k�������2{����ك�'v*--�>	Ȍ{[|Q�ゥ�k��eΓ���ѫ��)��_�N2�IF�"`����ڬ×@�&�P�.M�I������ϯ3��g��
�<yr���K诬���5�O�,�<��tO�t���:<�²p"�����d��_���5�������P�ǽ�-۱+���@/k?����ef�N��aʒE��B?ހ���p�2.�}	��|������Y�Qf�IK[z�]���9c��RI2�3�LO��t�2�l�y{9.�:0�ۧ����\�hu��\�f��C0���B�͸{��4M�	?��'��:�pKH��`��}V�����qeP?,Q�:��82lpd2�j��PG���hwkzY��t���W*�_�gG� �~H�,�%��,؏:	_ъq;�Rm�ҹ૘y��/�@��ʷ|��)*��y �čf�`�����Pd������Hm�n��fa�q�`�6640�=l��B���(����َ1Ј���&נ��襮�+��d��G�r�O�i��j���c���g��"/�1�&���I`�$}��M@�$��W�ޞV�����Ahv�Ζ73V�WEV$���]a߾0°�C9�9�m���Xw(�πg#]S��qX�cNn,�#NC��*J*����DΟ��T�xȶ'��'͡��]Pˋ�@��W ~^�R�m�aמ�� =�3𳍽�?��LlL2��B(agw&r��!�������ne*��nW�s���$�����ʱn)��E6[&���Y�BV�\}ٓN�?��Eb�-��^eg_�0��?���5���x�X�u_��g�g��BJx���D�/�Z�;Id!k�m��(����CCC=�&,�����o�W�߁�O5���$��m��mD�N=�g|����U����	|!=�O��wa�ٸp��ݻ���^G��;���M��a�N��sA���k���Q1�R�3�U ��fz�)��ZC��σ+������uu��R�1�t_Y̤-��i#��{���z{�˽׬ĳ'������g�+3<�}|z�����U�m*�S	���ѝ��{=��s�Nn�sh��e��U^���j��ۥ�ms�퇜ن^K�'(h���݇i�x�-%8c�W�w'���g�񜠟�F��bg�RȐ����c\��D�������u�E��b�[���3yWD�ʶ*h1pTf���`_���Z*�X�QZ�A[�zu��~�F6����+������u�T�$�\�
�p9$?O��{:��D.�+a�7�y���hpiz��d��o�Z��q
=�0F/�mۣ5KW���j����0/�������]���R�W�sk�M�茤DN�#���-'��� {��/��#'\H�3�;����R"Fϧ͆1���ޮچ��3`�z��F�/ԋ��`�R�3�����$ڛuf�e~�65���P`� �tXaaa�2*۱Q����x����r�7\?i��~;Û�gm���?���|�l�,�\�S�*��.���.�+�����>���F�����+/D>�7 ��w���؀�ʾr*���Tv5�~������h�
0$���$�i 64~�O7���Г������ҋ���	e��o�]SlS2�51-b�B�G<Pͪ��=�n#��Ed}ĈN��ό���ǡz��>觙����w��5�Z��\t� �<Ul2�Q��ɡAJ�"Lȅ����T��a��?�=]ݐ������?�JC\&���TVU���`a�;�����n��ː-����x�a4�fk�O��"
�Ӫ�O���a��huI�Xw׳�ޔ��|ZOp�"q���ҐL�X`S��+���;�\�{����i��n�j���AH�{h���Q|	屘S�����	H����o�nc7�gk#8w�W/F�����lڗwo�>oi8a�7ȭ�ϖ����(���~�Q�- X�����O�o`1�Vf@p�Ç�C�}��J|!ugH��81p���˫+$�������K_�S=}ګ����{Ĥ�U^����!>*t����u��Pob`*� �Ȅf�5��U��7�6��$�ͧ�P-��簧o@���	�����E���Y��
Z��IH���T��;��ҫ	��X�A�g7b�ïs���G�������X��I�p�!H	Yw/x��}7�����<���_� ������������A�0Ǧ�O�,!e�&�������ۗ��i�ii_Cؽ.�)�.\�ƺ�@h�����n1�_�����z���*�[z��({�i?���8�>E�S�m���[���/�8�?�����^��F�&+}��](R߾�<��gū?o��@�zu��nn��i�����3�R�s[[~L���E��U�!�5�E����V��x���/��V̲���j�}k!����kR���tC��������{���<]`��&�}۽3*K�;|u�C c_i�A�
}�?Hq�v<l
�Zf�	z�$ZU���8��0$�;���r�]X��u4k�~���LE>�_T/'���}��=�~9��+�ݻ��<������w�:�j�e��?as�C��,#��^^aaa�6Ч2=�!���.���v�[�Y�:��Ȯ�0�`wuu]�7}���8��)�P:�,�V5�/~&��2^��=�^y�0����(����Y+耇G{�Z�\����ϸ<�/@0+`��ݻ���%��>>>V��L ٸ�Cs��ѓ�kG���=�/��'ӛ�SC�1���37�a�ܤ��(���qWfG<��e�A��r��Ѿ�`��55�� Jr��?ɯ����]a�C���O�<���U��+ab����y�1�=� ��K�
QB��ʾ7�9��0H�1Ʈ��{�t��}��Bev5��=���Ð��7@�����3��UJ����h�ɓ`=���T���!�@O�q��2Į�x+ʒ��vh���{�t�VٗE{Iu���a&?8���H³���vz�sL�[����v���@�9P���)'�����*��@Gl\�������g������Q6�(��jo;�<�ﳖ~�i�����-&�xC�����K"�ǒX�����0X&a4�fEa�8Ӻ�����P:�������fF�<*q%���e��kO�A����Bʯ'�b�+�V����wumq�����pv�V���`�)�[�_~J\h�rr����7��j�m���n/����{��c!S��T��XT�ٰ�'cL�������$���돻��+R5[jV.���P�͘�?��-����ߕ���^��K�F��=�IiK)�G��I�����ݸ������lv��laz�e<K�T'v�1�󵥆,��eJ���tE��v\�i�!3���5�&��z��%���hU��a�С�y���z�3Ϯ� ���̗�����[�|��DEM���H��N�<x�F�}��tn���|�aӀ�P�����g#P����L�]�9e��4=�z6��zUK�2��T��e߾��i`�:�����Mv�"j�*ﺻ���ċ5�����/�)6���]�(fR=G�װ��O���͡DR��K�wi'}����S6���319�����:�莃N�u!�@�)�%��I����Y��#�����eΔ%��z�d�^�!h� gFLa��ֺ�Mfߙ����'nq�P!����>��ׯ�W 2��n�ėپK)-����E~����w�3��g1��g:�� ����Ø��;�Z�5���li6=��V�CyF�NUK�{Y8����Wۭ��ԓN&1���/�0��|��(����̉ҩ���މ��U���;����r!�1:_�θ����c���Y*fe_��[��#����L -&���TNR�] "��,.��'�"��4��f�PΣ7퉎��p2%N�������
c;S�E�����k/	'��wQ;p����b�}�yˆ�yyy��b�s��wi�)�y6}O�j�(C��aw3��L�bB��ڥ�x28�S�O@ �w��+ؽ�5$[G@'���-_�F$��"�#��v�(E���C���l6���B����&߲�5�p�`���o#�@G��m"'�����;�G����t��~w�2�Ō��ԎE�Mi��ω.��L��J���A��,��-�1��ۻa�ӄ�|麟`�K�)�W��˝��UDYs=�KG��XS��ڹ���r��J+��zM��F>��3�u��$j5*���.� c�����tC,0�&�j�28_?|�jt�1���%f�`�^�>hZ�fI{�V�.���t��}���c��]n��v'm(���$m����3�ؾ
>�v��8��s;��ʾK=@'(z�
�r��)�^�3��M����`�Z��F����@*8���>шE��$rnfĔH��$����C��-�g~�t��1eK׾K������(t̗v_NZj�垓.IXx�PV�(9�J���zP>�1e���TU
P}=�����%N�@�Y˗/����	�Y�� U���T&��\� fҘ�,rp��s��l�8��StҚ��Z��΁ ��HPbc��,����I��3<�@~��m�9�7WDc��.���ҧl�u!�l-�K7ٽ��j������{����Z����t�g�K)��/�Й��r�AМ"@�{�����C��D:����l�y��~�;�U���{�̕�i�f<'�go��xt����f�*c���bu/���rr���7�*U������/�VA�Z��V;��ɮ��-g+B�#_���S�ҕ����K/��:�n�H~���g���a$��
�/;����	ĉT�B2�+�F�b��\YY	5 6�\hs�9 ��gڒR)1�i7�)&r�(.̞"��w���w�v}o��&���R��m�s�r3ʦ�������Ŧ����|K;��ɟb�.�w��]��K�b�]?��CZ6�p�_olo�CC�p��q%��W};ʨx�_�Ź?��c�b��7y��5;5��@ۉ�*��gg�B�S��x�oϞ=�PǿC����ǟb�`�z�T
4g��G��V�$��Ӟ܆?��+˵��c��*�:'�wOp�z�;/�hS�U�R�H�bi�����_�� 6GOA�&-66��r}J]�r�a&��� ��[��WŦC�wy150�%�e�oy��^���"0;��ǹ!-/o0��f����7ؽoIJc�m4����e�%��C�hϐ-#+��Qh���.�.���՚.78_Cm�b��Ągm����Mo�z��'��ӽZ�:�=vlp߲uZ%{��Y���˽�� ��2���3?�Xf���'�f���~�ZDO�?�X/�p�gc��L�W�C����G'�!��Y e2@�HKX�cJ�t�����?���Jpy���.!�$�2b�����s�t!�����+�Ɇ��O��l��Z���9�:�3�v�RF�d�u���B�8ؾ�7��y��$ۛ��-�|U0��j]����DNF���	������l6j��@��=���+x.��,��-��s�.ġH������#0�z���DN�)z(�G�-��4�^g�i�ۨ�ϵ*�4����ad�B�E�̧K�<�\C~���v�W�!�L��E���JA����FV������|l}��!�. �� �)@Ȉ�nu�y��[]�����(^:[W�U��, .��J�֭�2y�������mG$$���z��W;��\.5{�@Q|�)vRUU��#d�;�v�o���Z<]).�z�=�iE��dݫ#p4�e<ߋ`d������:`���l1𘩓��'Nt��5��>755�(��e �(�����#s$�$��m�Q~�V���葾�~�������y�xv��SF�����z��>��C�8#�P�p�p�o�}����P;�C%��Փ�i�����p[wh����𿘙��[!D��4�k�J瞷�$�]���X��#�^E���ep�[�G=б�!�I���e.$����ci������qM]������^̵*�ԆVM��2
�F��AAA N 2��`�%VD�j1�̊�(T0T�APA�L"��[������__�O�9���zֳ�����L�Y���SxO��ZN���G��N
��	^|�<pJ��3�۠�����ň��^��#�I,CP��LM�/��+�?����G��/�?0� .�XV�dh|2�����������Gث��|=yZɧ֫ҳL&��!0��2cu����*m�f����]�;�&s����:g *s���#g�m�S:�u��0�\�}�}x��4'���a�.��'lN���a�)�����V�Ovʔ��t�w�		�_��`z[Ҍ[�!��� #Kx0�\��0}EZ߅O� ��M��\��Cx�ds��g_G�Si�A*�����*�'�r��[wr�e�]�P<�^43p�,`�d����pM��%�kT�[ �?���.an�.XH\�A�{�+��qƧ����a|z�E06;!�Z��͵j��P^���������@�k}��u�?�Mc��5��|�i�Bړ�>|%<6[�I��	�5��M,0Qe�?��7�X�]Ӕ���1+ZA��6T�zt�ᙐ��Q�e)��N��m����`v���'!��	��ط)#���7 X�9g>��T��^O� F�wM�*kP:c�-�����݀������ܷ�&�T����\��I&���Q� -�Ak�+f|W�`�ҥ�8���I����9���3�;���^S~FY�f�1≚���d���9����`S'���գ�F�^4k�����N���egAޔn���1>J^q�l+K��b-]�l@S9 �bA�A��O$�]�<b�!|Cʚ�k�8%gL0Xq��7��
,>�=y�#&&fҜ�����eK��ZY寠? p����cת���]��X��i��#�v���6�50�p0p�f�P�l���~|euO#�9�H��Z���^[�	��o�+f���>9^uZ1V�������C��5檧8��z��ΝS�O�'߇C��%W����6�u͚�oͳFSp�!�����9���]�-zwx�MjZ�h9�tXW���o4n���U��w��T����������Xw4@I�%W�*j�r+�ȣ��°Z�^��L������G(b7�KB�2^W�{�tԷ�F�_�����GQ�[�����������v�j�{M�����u�=��uO��������{Q/���N�_�����u���_�����u��Y����C��#{����3rW���O���[����9�/��|as���6,?j���Yk�˲ϼ��t��DZ�W����#bΆϾ��U��ϯ��f�E�/By���	�w88dH'��9�p��`k�Le�}�k�@Q�ę���_����_�3��_SX�o�,���O�k�B�Ǧ��6��V��ٶ�m��L]����6�?�[�M����{�%�s@�V)���ӧ���F����&���@Ly~�j�@8׬'ۘ>.�5}#�����~GG���/�����gI��>#�L�m@8}�}OF�	+���z���bt�x(F���Ƨ׹̼�}=*�,tي�ɁL�ŏ�5�o���~�F��ܿ������
4���v9���ٷ�9�'�!��ۙn��^�~mpgDZd`d��?���eJ��ۗD�Oh{���̲�?V![2�S�Ϡep�N�8*�y�T�g�jGo��CP������?"!�K���1�C�a��9t��q��Do��ϣ��Gu��{�4Ķ0�\�ċM����yh��r\>v���hF�#@D�h����T��飀�tS$=��`��:8U�]��!����8�}�ԌN�8�?kkk��r�lf^��Ũ|�/�b�X�)��	1���z�s��?ߨ�1��ֹ���wCv#����_D+tF�������,O�����F�Ou^����*�az�9E\�%'�3�����������p��1@��󁱉j���%<$�+�Ģ�2���D+�$*�dg��V4�[�'�4������G����B��#�4g���֧8����7�j
+R�v�iM醴3�G�	�K�� ��KP����$T3��j�;��v�n����	)�4n":M�'��Fʺ�j.�A�^�}�1��{�{�/��ّ�D��+�^��$��>���l�x]��M&a⍏v�Lt��X8uK~&1����j�i�Lm.l�P���,���MnC+s>=�6>l�ԝY�R�kg���������Ւqg����(�
^s����l�d�����)f��Q�&�i��܏�8��B-J2J��-���)�d��~��=��u���������og������:6{�w��_��t�Z��i4	w\ł��3O������3Sګ���簟d?U�
N�̑���9:	"2�p�!�$O�.��?t�a�^lT��/d�w؄Y��r���ﮮ�Z�?���E/~�P�p^�����|7��޾5c����B	�՜`w�

F�9�3+��L��|��8u���Q��}��FLY���j�1�"b��T�&;%���fP�7g:"d5=C:|�O3?�j*��Mѿ�iuR���$gg��g-=VR��4j_��-�90���~n�!��˳��݄�3����gI��"�:[pz{�r����jbc�S|9��B�hyh�դ��7���8O"y�}���h.۬ƺ���PxA�
&�o؃��P�6�b�!F�h��#.e֎�
��c��a"n50c���Z�i���+�٫h'D�7Ϊ�o�q�����Iw�ol k6���>�-x�&��{H#���w��3c�W��&�$}ô�A[[�DY��n�g/Nu�}`}��Eiiig*��Q,T��p�#�L���P��V�w#Ć�j���-�No�J͍y������^q�_��c���4Id�,Y�P���6]ʲ���k�k�.�B�/GsV���Y��Y�C7� ��wk�b\C�A�|�f'纎]3}|�Z����>e���DEB�O;M�5����a��}z��2���g�w�Đ|�L���[Mn��c	�t���4OO@ZZu��0�:b�'�~���-ɹ�a�+�b��\#����n*�yH�ۦ��/f=�p�/`<�|5iAX�ʹ�G��p"x��a)|p=wy��]���bܣ`�`xnH��N2�� Y��y���[���ʇ3d�XK+������	���^�jFo�1�e�����$N�
8���Yk�U�S�Qa%�t��8�B
>��S:D���#���#d/��Z�^���P^O�za�(�{!���g.s�7+��9�����#?�b'��ь����_(�ܻ��Nኸ�S|yPik�8'���x���J%C���rkW���|I���3��s�U�_F�17k���1sV�8i��T'��!��|\�.)V��f�b�Q�����o�ˮ�9�ai6�z��	�BU����}���`��%9Df_��ڷCz��7���w2���8�6�Uw�[L;�b-�����G�v4U��)@�v�H�)�u�J�_��|��X7s��d�U�ܚ{��ߐ��"�Z�w�054ue��_��u��]�>$IE����� �'�u,��*�:3�QK �^b�[�\��VB"~���f���r[[��*�_�[�]"N��FB���gM��0��A�����3^���gn��Ө�Z��"<y=��KM.d+8Qx���������i�$S��<�h�����a���<��x",1A�3��R�I���*�i?���dTjn�^!j���}0'��?������<x�WC����2������bG�k�J���C��Ei�ָ�L[���;��Y0���� V*1�j�F;�-��Էu�t�K��N=&+�M�)�W�;�޾}��G9�C��kLdZKMp���*~�:�1Q� �f�4��n.��c��%!����B�_:g�ϗ�qvd���� ��Q��Ʃ<Zql�u��9�!�����Z����<��
@���W���(�v���@7�~Q[�"�6y�6+�WNu͚�M�h��jxC��3�J��Sd�����(��P;ԭ.���� g������h�&�f�B 6A���]�<]ݨ3���y=q��׉6U�th}K=����Y]Cc�d$��n��}|��I�a�o��!�h4�	���0i(kE;cx�.�,�1Hz�Co�x����F���K��P�e�XU��sTQ��c������ȼ��/Uh} P�wL��,Y}��9�\Ń��)<Ip����}��	�ǻ\��2Ku�=ň�U��N�
a���~��S|hnm,"v������M8�L�I�h�{J�Jg$/ԟ�"V�k���w2�b']0-�)W��Fʚ�;�#'5:���s�Q�?��E��a�l~� �4c�-��w;(�%e���%�����N�"˨�C���⫵ַ���$��bMM��4����i7�$���0���tĂ�!��p�,(����zP03d6��Kq�r-*gq����O�T"я"��'��G�3Y<�p�ѽM���G�������xʑ]>�M�S��s.�*�`�� f�8�����s��K���c�qIMv
˯-����-�`dT�`���i��qf��\��:�����Mv�oP!Ϭ}gblH򱍢���^������'N|�2&�l&Q�=���>�����@ď�ZC��#�6W��3�(�n-��i�&6%�*�<t�o_A�@���U�O9�s�]""�VN�T)��2vtu]��{oR�w��^]c=�F��5����D����	TD�i?�%��c�
�!	�s
��7��QN��Du���9�c5�	ze�DX�@��4�J�����/���ǂ�e��+�h��{�nH�]B�.�	�_�7F��{f]ч*�T����(x�~{���sY�,u�TU���Axa��֪?-�*��P.������p|�wASwa&�t�������b��:�@�d㔗=�!+v��O��}uGɔ��l���9�0!��P��Ԏ��g��V��Y�{��r�o^�EW�M�D3�`��$���j����.Ĳ?y8:B!�V"r#"�����["��O�c�yT�έ��C#����"�+h�-�|>�d�o����}���]3j�#`�8!��<�������0B�o�V��C3�Z_0�z~�bH�d�� ���t�"�@0��숏-S�G��
�����1���������E�� �����і��~��y෥-�Z�!V�&�3���~J��3c��h�S�D2��u�Ʃ�^����r5�"�~",|?�z���������F��+kk�Qf��
gx ��Z$BLk�f%��AE�7r����pK�����_A�|4�����i�|#�_����U��me�� ��œ5�!h~\+`��Y�޼t�&�*�Ar�Ko�<��ӷ�I>"�r��$�av$�@���zF[�a�ϲ���V���n��dR;����d����Ċ�;���둟?��"ze!�-ʭ��G�����]C�Td��Oj}��k���ca�Ȩ�ѵ��jA�P���P�ݗD#�
�E�f��j'�@&�Xx�j��dV�K̜C]��b�!]%I�I�25��k@�����i��z"Bn��+Л��Bn���y�������y�xǬ�F�$l,w"l��f�[x.�gcu`�[DKA}=����}��G������No;�)���P��n쨡΅Fhmw䊻�W���Z�Fn��h�e�DrG?���{1z���s��ju�3�=�s�A��Nar�j�l�x.8���ܺ�����b�B��#
�O^�׶���Y��Y�<p�`<U�vD� m=R��+pwV]�ۇ�T�@|�)��"����;}��i�8Y��? IMI��n���H*ѹE�G*��=C];z�Nސ೤>��N�u�uV%�W�0^�U�{�5�.8�t�j���UU�=�@w&�<γb~��w��od	��V�w��]�J�������ϝ�1 =9��\��7C��{��
��{3"�[<S*Hĩ����k��)j��c˱��щIEZ�M �Y��湘D2Plp9|��'���MU0��O�,p�W��'��u�A�!�Ԓ�7�����.�J2y$?��ƶxnm�L���\ L�~z�Ed��()��*�VY�K���z�����tp����<ȳ�`�q�ݖ<�!������O�U*�&<C��5J<�mV�Crh�vH=a�z��/p�x��|Eb�I��T��ص�Z3���8�����F>���=6.����f��:��z�ʩ���"׹�)��i!)&�q{"���mn�ھn*ֵ��O W,sx��6Br=������9t�C�)8&4e�k\2����(:\0��LAc���]�y� ��?��"�c��0r+�8\�F�A �v����
/����*�s�U
W���B��P�*���$B �d�������I����,��4���])@��vT�r��j�>�Ľ�$AEc'�Z�㼿����[�G��+<�]:68H�S�&����3����x�uEv=��0��1�F�'��k:}2Oq6`��=�n�D��Y٠LQҳ6���h:Uk��� u��x�D{�;���!��"�j�&\������ys�ۏ����'�e��Z�z�d��<�B�6q 5�������{�=�}�<y��zx�gQ�S|�9�[Šy�3+��}<;��J`!\��O���:��~�4�xH��\ױ��)�����F�#)�r��AF�}*�L�mOz���dZ�\o����w:gdQ�r|��ߞ\�x�%��+�@wCe�񸭭-���R�"���D�����v���V��D�s�����V�����C��V�������Ldޚz�!C���Z}�9�d!�{�����u�{ċ=�E� 8���jU��><�ם�~�$;����[B89u����R�%7����@��[*��2�������ތ\u��ӰЙG�Y� =��*
��_@o &X��oW��^k�k1��$�P��`z����d�L#��6�+�e��`��A��Xj��k	6���w7NQG|�\�����J��N@@����N�Z �a��G5d0�r�V��.l?t4���¦&�d����� &�b�	�`@�?���H��df��c;�(��9e��U�񣀂^Y]�- �JT��v4��խ�2�J�GE� <��{X/���/����f��Pu�ʅ�"k�2��MS�.�!(�ؽd�'d��'L3��vѥ[���+�	\OR�#�Y8�y��.�707Ћ��%��y�a�������U���B.�1�ălpd�
�v�e��5kB��IO5�؇w�r�h�~��)،9� N��9�1�8Y��.j#<��
��^�$jI�hy?����c�����b	� i������v����R���1�����T���f���rj�\�_��	̤;�D���Ŀ��7�A��1a�.��呉�"h���9w=��f���[��ڃ#{���]�KcM3Or���Z�#�]~4��ٮHR¯F0�b��L?‷��˝3,��	�%���i��*)UN͝ĥd����θﳳۃ�ɓ��U�;���ڿ�H��x]C��{B4<����%n�@��%jo�ZC-p��S�d�纊j���Yſ�G'�ן��T�*Ů�CWV����g��˷Я��~���7��&͙˔��'*G3�?��Ƹ�6gg�&�j#K�2Y�qF���%Ү�Y��cܰ
�1�b�H������j�$�n�eȟ,�� ����<��c��j��Wϭ+�Δ�m2�ـb�ɻ��ʓLNr�Ѻ�;�@q�|�rZV%�����ԏ��ķ|�����#�q�b�G�fL9zz��R�qC�J%���x�9�<-k��9�xj�	yz�59��������x&%����m�_���ᾮ�ݭ�X�f�uʻ�_�\��u�$�rv�Y��	�-��h%�h�(sӟ���i���2K�:�v�.j����S���*�}�\����]�`}n-)��i�Dm�uW��2pΘ:VyK����.���p}(o��>��~"��j+�]��V�-����
�/�:}6=�H�Cxƀ/��Y�GUH$Y�eN)	~����{�>]���x0�G�7+hy]ӑ�/s�Tf;�Q7(G �R��X��$�#N�-@?{��������"v`���@���1��V������  ����!���X�.j�8\%Q�?gJ�t;o|�r︬^Ї7������V�<��K��g�xj��k���~�X�����A����f�5k�4.�U�M�M�Gt��BH�޸�+�HĂ����z���he&��(���O;A^�m�99@z8�vБtʁ��"哜)��\�MYZ� ��&����Ӳۉ���0^1��N<����d�J�&վ�CT\��fB��;)���v���ƣ��4�P��.�F���^kk��eȈ5JoJ6��.`��;��ς��gΓw>��N9g�Ds�!%��Zgrgh�x��6��tz�;-��0Km�� �έ]�r_<K�2�����z��Tq4��"�=R�&�k�{&#=]w��G���q4㰚���ŭv��u]ح����D�d�P@(.���#��c�tkl/;�Í����OwU\-��
0�Δ��ǳ ٝ"�M4n���Û7x#�B�9��궓�
�ҡ1{�S���ܹ��i�=YH�]̭����t�lěR��>��A�X�b�8��S��z����窐���ɿ����ɝxg���_U�rJ�f��<W�|n2��ޑL	.�O���B�qq��x�]a�=��$��;i}�fL���r[�̾x4C)C�^;�6�CPQ����P�䆡�7�lw��(Gs%�+KR>�A���j���;�K�6݅AE��4 ��|v7�6�;�1^�4^��MA�f����C��!f��!N}�ZK�Z?g�Οs�'�R<Kxw4ws��e*��<wI$�Q����1���,����/���e"ea�ki7����9c.� ];T~U��.?I��S���p�52
�E���X���u��$��5�hdA��zn�n�5�� \��oBւ{O��cG2.����Z�F�P��[;�{)��n/�*p��3�5kV�Wz�q,�ꐦ#ꣿ0C��eg�3 Fʔ�z��.)v.]u	�H4m�����)\��L�e��kޤ0Vjl�.�tP��ϭdq�,�@��:��̬�o�،Z�B'/6��o�d��*j�ExqwT�(��v��S����oS��t�ώgJC�&���<w�������'�SsuW�d�v���{�NV��$�Ҵ�u�0�D�����n�~��7ߜ�|��W��׮s�V�}I������;L��şUM�S��_�L�^~�T3t�[�Hta"�,$!�5����*�ٹ�Ф�F�Mj|C��:����&"n�5��L��I�=8���|0N񶅄�x�/a�@:�x|��]�i�u����$(�R�H|����J�C�8�Fsd���Z`����T���d��`�;Y��999�H�l�,P�F|(nz�X�������D�B-�����V�)Y|�R7�?�y����G�h�Q R���,�K�#] 2]W)�����M���
���C'���+�DS_�b)D^��l����K�ńy�D��Ժ�7Jػ��Y@8�gu��<+��
�
r�;�-:I���S�{���lv
�*��������IN���"�h�irйy�I[��'�.�j��`��� �H24�M���i�G2�O�mm����zۭ����)�D��D����be�:��!��/�tr���e�q1hi֍Ρ1�Xr(�s4�9�0�N�8�O_���Q�d' � |%�THMgM�;��������$i�������g>��6Y��� ����1� ��}���aV���aU����� �'���^)���E�˅3�S͂�´T�\�y~��-�م��;��Z{�E���bKZ_%��d/��%���Ǹ2�ءx�<�u���o@oS"?�J}lހMW�ˣ�EZ�\0�����r�!G C�*�b�H����5/\���j��&��	*V��U��N6Z��!M%��s�����po#�������dtEq��%���]�5}�'U㊽��y���U��c��'9���Bh��>���L��M��;�����@�.�(����L�;{ɚu������jq�.��z�����o�tU��8@��ƍ�Y��T�GԵK|H޷�m^��#��f��ڙ��ښ_(��H�//C���Ul��s���!��Yu�Ν�)V;�$\�%R^�O䚺;8�7�q[ᷪ���N�:B��<;���_싻b��ڨ�k�OsTH�}x�숏�m��Z�Z~4��Xz[)�s���c��#���TT:?��+�b/��j��Xs�G&q���5�xީ҂�Z%�]f&��/k�@��I���-����nV�Q�MF��!��pwM�����t���xyc�P�+��<�l�~EQ�/D�c�9x�,ΰ�m�� [T�-����� ��l+�'���������*u��8�9�L����i8v��	/� ����<��LwK|;*J<�Y[ʭĦe;axF�w=���g�ٛ N<~C\�V�V����ż�D(�KX�t�J��cN�]����U���Z��`\��h��:�9��h�x�~������� U��Vnbbb�An~������g�7�����v��j��0�#� YWSH�M���c��FDmOҷ����6\@��AF�P�V�����/^�q��mUc��v�$}Y��v��� �a�U��Se��Ж��*9�	�!���x�椦Ǜ�%Gνȭ�d����jr�҇�T��p:�kc�U|���f���9�=y��"�*�U�35����-q��D����Q/X�1.A;��F�*O����x$�_���@�^��VT��.3��p�%����XyC���!����C.ZN�ws��a�O��8W�Ɋ���F�vQ��X��Z��B����{�/�����Bw�.#�_��W���#V7v�*�\qύ�ŏD��0�^L�����4���3^W�W�C�n�iE����"�\�;��"1���N0s����N��ր"�בU�PQ:�s�#�1W�>������ș̉"��u�PO@�0�6v��t�N��DsE�l-�w�F)�[�� �I��At��9q��ض�������py��dMN�^��^�u�P���Tr�1��ł�Ps�jHDrx�@Z�VؕR}G���:��!ƻ�/IO����16nN*mgH�ۈFoذA�!׹����;�?�7\&%��8�ܵ�5��rv���IM�n��l/�^�n��y����m�B-v�!'YE�E#�&�;��hM]��b��J ���J�"n֍�?n4o޼3�?۲gaX���Γ,����=��t7�ߙ��m����0Ƿ"fm��a�n���s�(�����n�� z<5�fEԬ�����$�a�ؑ0t�睇���(�ޮ|$�}�nU���V�/�懲?=��v��KD��Yuc���ywA-fB�aI<�x���xf�r�E�1�r`��7�\���1Ѐ���ܡ,��������+铹��F�����M0S� �\�~_[�5!����3_AzLK=J�?�r||\bP����(��c.v[[��������4^�*Wa���]{JC	�K�
��m�A�x��Q��t��t�q�DE# �� |
�O�D�,��q���go�<I�w�~Gw[>������%��)��c<�S��U����P>���J�i�%f�Z��j�h9��Wɟ�{!�Z��^��~���۷�3�RH�W%s�Ƥz)>_����ꋂ�6;:8�-���Ӷ���r_M����Էo��91��N3��9(m��s��~�Y?kE#[-�C��
zX�.���Kz$�H�Q�ACc������<m��7�?�$�1�qBU��]��)U��\c[Y8ىsIЫ5�����a���4���q��=6_D�Ưt^�O< :�3�I�~�o^-E�\0�3N���:��g����C��[^�^Iv�[NS����\�≰�����=CS��oI�	oܸ!��#`;�D�Wz�)h}�s���f�"H���ma�����nM����e�G�Պ�����N��.JN^�)��d.*Q�����FFE��nkq��)׸�~c[���פ]!��2��>3&��=C��(��C!�b��B�]Hc�o�8��LK�_�8[��.��c3��- --~x��Gu���}���0m�~}I�}��m9��#X� ��B�Ēl}Y�����r&��	��Aa�5HA�C-����R\剀�*ȃ�֛�T�ќ1|(��:�GmW17��^:�v���n��8��v�T߿_�W�{��.��,O���ػq]\BB�����,I��f3�-^�t�o�D���;xh&E��qT'Զ�������Ҩܮ�;�{z�.@_�s�l�X�ds�q��Jm�ۂf�ޖ{C�y���\S�=~%$��:�#>�Wo��8K�1בCK������=��`.�ؿ�!y��ɑ*\������}p_�i/������E
���$7_�9Lʄ�9N��X+�J��+���or�;��_�/X��R����;&@�Ǐ�l�	�\�!M�$��������kM��ڎf#V�-�t���& 
�X����*A����r�o��/�~5eO	��%��~N�^t����?�=ͨ�w�;̒�#_n�H�Ы�J	���$Y��\��P�ot�e�|)�e�A%�*N�&��u4��X�5�r��Ns�$ �8��l���F������e_xu�Cu��2���[d�-��{��"�d�=XQY9�t�"�ce2��	��=�~�+�t){1���z�6�4�2GDav��g��
�t�"��"Z�q�E�]����=�ooÀ������&�_]]2�F~�!��#��A&�願�t�z�h=ѫ�{3f꟠�Z��9(�"��jf�'py�#.����;B�������|F<h�jHC�:��%=�� ��=��*�~�@��5�:�V�d����T"�[��EP-�詝�{8��<(�i�('�Y,'���`�N�e�e>�?ϔ����߭H�*a)7��������{�lU`%�����/�o����gn�q���N8f"���'9yP�Y[=���y�\��A/�;l/���8Smg�k��3.쉷CcP��X�S��_�z#��E�/4�͊���TX���խu��Σ6W�� i~��+"@c9C�a��H������RS���t�'��IMN�G}y�״3kp�馬�.��k�LSn��}派>Ҁ��@(Z���J���'��;��S@�/���@��o�x:�y�9����qz/{�@��>���js5��:!ۘ���<���D�88:�R�p�@�uy1��Q�zL�C~�%aw!���-2��'kiЛ)����Ց����A���`��V��-�M�՝!P�w@-��/ߏ�	�&$�U�Vvu�4v����~4꾽l%2�B����J�w0����Z���}��+Q�M_+�]��N��XBs����䔔��4{���d/Q��x���T�Y���~�ǽ/������m70x��U��?��_��B��X��X9�� �yy����)
%����n��U�V��*v�����GF��݂���'&�E�L�jA�^0�nL�'�B0h� �5g.҈�O�AEy���޾}{=��k�z�k|{Z�P�E��7����VLN�eյk]��K�LJM}��~f#��o�6<���'���Y��Q����b��m�k2�����S�R�l�d��ոR�޲n�b0JB8�%[n��'�����ݬ���p[m�b�466�T9�+~��Λ�nlvB��\��"��b3��-�u��+����׵ҁ^��_�iu<i���ʉ(h���?��K v��V/+;�#gP d]���Mv~�;�]<hj@��2��'�F������^��+���)�o���ɉLNNN\F�����m���>.�>�@��\0�x��I��ms1y���)��	�͖T2�Ġ�$�ۓ>��w����F�m��p8�ug���`��㢘����?�DJV�dL��Z��V�%.5X͑}�%�����<�
�b�r`u������5461����TI�8���\㐢օtV5��oJ�t���~`+�ң�/k��5e�=K͎�N4��73$�)�xb�#�V�̤��ο�߿��x�|p�rՑN�St���������Q�8ȼ��)M��rcN�� ���.m
��v���;;�����UPwO��M;�%��\ӆ�O�)5�� ����(	�f��]�Ψ�����t���"�$�m�*��0'Ȩ��d��-��S��<Ez�{�9��;B�J$���k`zauDQ�S4򕙙��]H�ߒ� �\𢳅X����"e�3����A�Ԣ1��Њ��T������|x�l�QuH88�x5}��!�����-F�A���MTX=�!�+�U9��]��>l��=-8O���휍�~Ƞ�5�s�H�n?��<�D���}�)��n��#�pI����P��ӖF�/ ���Jt�])S�}�$�����V��Oq���Y��W���>>W�X�.B���[����jH�)&&Ft�#C6N���Sk^���U�+�ַ�n�}w����r����c�'�,s��L�Q�JM�^��;B�s$�g#
']�4�=ڹ$����۶�~	��Kw���$A���O�,m��C�C}(��Q�&��8�<���(�^�����f��5Kg��`�C!�Z�`ℍ�7į�!���"@1��5��c�菺C��L��NA�z9�3���e`ʪ���0�F��e[|*�7e�*6�g�M7�n�V�
��C��E)N��\���2kf��x��f:�3:�
ݍ�X/�O��>�-�ߏ�톊c	��$�m����J����2h���S��8û�+�w����^6�N����������r�V�aS16n���^R+X0�р��X������pR�_<�37��{��ؔ�Cv}����fnn�������~	1kf�MD�>��z�n����\yЀ�m�kÇc����s���R�$��Z�
�>���Fг�!}�h�h�d�\^� ٩����x��� 6,Y���W�LY�f�_i�;B���=44�CY��1�-LY�'�R��ݝ.���D��{��x�2uo����e�@�Gjq�ũ�!��9��sԬ�0��� �w��߀�2uqEG�b1�:�b������"M��)6���U�`Zp�X�f�o @Y���`ƒ�F��׼,�}��Q)�F����~/�e2���	�V��΍�:��*�`�%�9�$!��ipJ��q1��X���a^�񃤏�$��T�����a�ޛ��BD#�8q?��LJ�UՕzc����u��aFo�!���f(�� ��s�tv=��K��R���0ώ3b��
�ߐz@���G.���o��۰"T\倫�x�+����;��!�?x���W$H�Ɣ�	�h�ş�|��r�dT�p�������*��t�������]ςҤ�������HWl|�/1�h����省5���$@��F́%oQ嘰o��u������w|ZQ ��ݘ��L���n���+��p�S�w��0��	�~��-���ǕF��O�IB����'�L�^MN��s?nUD,� �����n�h�0^Oc� 4X]G�?tTi{̭ʋ%-���9G��K0m�G��D��2}��w>�u��c������q�{��	9Vq}�Ob���h�X��1P�=yv�C�w�<�]�o/)�q���	w�F#o7��Z�ͫ�!���a�ޥK� ���/]*�����4�#Ô�;���Vۿ♉K���ݚ<yf�h$��JM��6�������&o��9�l6P�2>v�Ҽ�[-`�(����R�̪��x��O����=����\������-r�e��Z%װ���Z=Rh.���O/��z$�^�:ĂP3�?���[m��`%�ǜ����ً1�nE��N�9Jk36����8�/I���ua����n����x��3��i�[�����w���Sg���eY��T�:\#��f��T��t�������epc��wx�����^�E�a�<���nk)=ʽ	�$�l���K$��20(�X��5���8 ���;J���y��,�^������x�,�K��q��Kc.L]-��%d��v�['k�E��c:����Gg�wے���T�s-o?-��"�+7�sT��U*p���Q6���-Ȭd1li��]�X�iZ)P�'���OU��\�ձԀ�W�Ph)y9o�<��Po�K~�k��3�#(u�4�(���$��	 ̖֗���?q�>ڱu�E|�/�^�W^����:�k
4�K���L��.��:>��a� �S�U�f6\7ۼ%$�v�k)R��o��R�Ӆ���P#(���T����k�<~�N���<@��n����oܪL�<�U�M���z/�6�i����[���Iv�c~8�?
K#�x��jP߰��gx{����ʵdc�ص6��:	���	Bh�+KG�0Gr�8�8_*T��z�^��Ơl:�{ֻ� ��8�$����ԁ��@$�ƿ�O`s[[�XZ�v�nL�ݩ.�6*,�r�����MI�k�t���ľ�>9b�p�����n�C3�̂�_�uCA*���>�L�YVJ��P�:�b�4G����1c�Ds�M�]�4���V�N�k�;�����b;�nvb�@�rlb��Ǘ	��%��ذ�n�yvħ2D����g�T�/�'=�a��U�~b��FL�1T`�&��L�{�J���4%w�M@�<8Lg!�fT����	dVpI�@�NL^�&�ZAXIx �M� �����OZ��2���J[��(R��nO��\��E7�E�l�c�̲T�����MS �?8uL'��׶Ҡ�O[������P�C�O'��*���'Z䡎Uo���� ��j��?t��_���`��S�^aSw�ǹ���=���K��d/�T�S|kD��t�H��)��dS-��xb9�4�����hn��d,�h돈ke����V�X����:\c,��73:��p�Ns4� dt�J]�P����EH�&�ŋM�w���`�灻�WZ��u|n��˨�׼�<�w�o�^�>���%W�� V��(���V�me�rx���+ў��"Z�]_�:�dmo1����ԥ��H��y�5P{��l���(V���$(�|,�*��k���;w�4d�ޚIJ%
� $�4H2���m�Z����>G"ض8���>=����ZD{�j�f̡��A\_�.���` ��p�~_�p��+�䒝#p��o���?Қ2d� �nٯ���g��� ���\~����[MYueǩ	ͅʮ��7Kȡ /��Μ�T��X��*T�u=�Ec� [d���t���O�6D�R�ee���GP�0f���1�.'g��CS�dk)P�j4J�*3HUӛ��'������r����>���CJ��D9�=�����L��s������A��vˁ��P���@}����I^���7�]�8��q�{"��	�����L:E�m���Ŝ|j���@1cI���50��^q���E�~aL�U�� ��ч�����L�ڲ_à� D��tdY}��w^�z[-�*�SI�4Jmv���ߜŃuޢ�yY�D�j;OY,��L5����'�����h�#}~���W7ꯂ�~��s�+�:��a�XH��U��m F���$�w�����Vi���[2�m���E��-n�V�sAW7uΆ8�b�eQpQsʴ�ӑ'9����d�Y��슫����R���k�9���{�Jp?��mn��J�<w�U;����r�v��!����=���=��ˣ��Sb��X�S�ّ�6���|�Q�z�WXr�;�I��l�	�0SZgn~Xeޢǧ��`B�+������p����E����i۽�"�)at��1_��|>��&�ż=�A�h���V��������~��W1���㏏���ԡK֓
׸����k�S�M�)(���Rv/m�,#۳����DRr�bt��ۡ���,��qݘhS� ���7�ꂨJ$��Ad��c��waԠ~I��&
*���fN��/�$p',ڻ@{Cܟ�r֗9�k��X���:iQ�t�߽+�і"��-��պ������)���t��"5�Q�Z���?�i���F�����{^�����}��`��"��
ܖ����J��W�qW���I��"z�N�s�AϡH��A`n\&Tq�h*�-�ɢ�P����A�}AS>�+�.xs8}1�"�m���R�̢x#�`Q��d�VG�J�,d�3b{���U�<O�yeT�,b�it���%K��|��}
F��f͚�.7}R2˩��k4V��h�W�50�|x|`~���d����Q1��F�)��9�C5�@iU�~W�ǯd*/�)��S�}���-yQد����{�r����g�mj]������w۷��Ѕ-[~��}�p��rqפc��������t7�<v����f��g׾����z��eI߰Κo�f󎸋���-{b�:��v��M�Z�T�6�w��0saa�b��]�y�tȘ��A-�L&rh��g!�p��Qn��	��A7F�U��K4BI~Q,�B]��J �_=�����C�]r��t�*�����g/�,�/r���Ц?����o��%C�*�]2*g���i�I��0��c��Z@�<�f��%�]�=���:mᑨ�o��[��\&���*�����v�W�Gs��G��"���Ȥ�T�|����"Lt����� ���%����%FI��l�o�v��������������������>��!��b�����agJ��5()p��V��z����r�����%��	��F@?1dund!Z�O@�?y���'rh��7O�h�0����=Β?ֺ6=��V-n�<�X��zkv�5�����f,U2��/��E~o�|��� /��A�`��:�ABf���?���bwu����򿷠R8���MSuz�6o��<�� #�ȝ�m)�(謁N �?���FP�p�&a��<-�AW��Ha8��!5�w��dqw��'S�j��cZ2�_�z�����Qm���AO� [����V�6d�qe�~fx�A!�u����=�^���䋹�u��0�"��KHm9�!6'�[9�{�kVOg�����^s�a}�X� o��<��	L��ߎ\��;��/�J��B�@e�9
�����T���9�Q���x���Om�Z�0���
4��Oos���I���F��G���懭�Ofa��o�>������l�)�T�Բ_H;OE���--�4���y�{cB��;��ޣC�[����w #j��{o����_KmE0���l-�b�*����FdqE���Z%nP5�b -*�"�5��!(� ��Ⱦ�gn�������>|�sg��Y~�3g�j�,U�G؈��2KJ\�I�����$
љ�|/d��6��p���A���_��=g�d�/	��{�S��e��K���P5���.��y���B�<G�!�LL���?0��hn�2l���zp�ҧ#X��XZ�͔�at���,s����оw7����%�l�@Ǜ����T�|8�\�����Iiim�d/���l�`�ue��D�YJ�<�eXQ�
�zs�����庽�]�U�y�"h��uIOQ_"`R4�	���@����.+Ds��~s1�M�C�l�I��V�r�&���'�a��z5(i�����W'^5a�^E�*hm�����z( <P�.�S��� �% SI���[+���3_ �}B����ǫ�7N*�w������|��M���~*U�BLXM0��
�o�A�y>�%R�v� �4��o�Bz�?�key����%�d�!J�\�,�PQF t�3�R�ͮqz�a$.�|���C�LA��W~��·�U�0�bsʎ�
���t�(�#�3�f�?�#wN�L���p��e���ެ�7S��A��?G��_X����t˛������Ouva����{�6�����49�����ZA�tǷ�ѹ��C�/��� �Ff�J���+9EQsxW�e5T��<��Z'Z�Y����O&��-�B�&h8���U�Z
��",�)`��U�
_�����`�(Q��5�xK����� ��������c*p�]B�ښ�|��)����|n�Û�s筟$����u6ࡗȜ*Κ�?��'f���%�*�����d+\4N;���k�y��@�9�"��\y�M�����!�Fk*�������>xJ�Oy��MA�'����6��#JO���D��dڶ{8�B�P��BC��iI)JK[����;~���Fi���$���5�?`�z��FZ�%Nq @����	
c�H�+����$������-kT�V_G�w�D@cJ�_�	� ���C\CŞ;f*�@����������%�a��G��źl�tj�OJZ杏�6y�,�`��Ot�h�ӿ@�z�ӭw��J���M�t\�<��V_4�/�HSY�3ԊTz��,~�h��iY�8�����5W�f�旹�-�v���]� �cG��N�e��1�Q���u�FDdJ��s)�i44� yd�4^�}�ě0b�
:IR�R��p<K�҂Ȍ�EDZ�i��:Y��ƺ'�
G�����]�L��p�kx����T3�����	���xV�ۙa5���#ګ[�a9����~��I���o��p[�ۙ��;��[s�j�DK�����i#d��`[�C��\I���
��Du����1��е�)�[91�]��cNE�����~�����%z��j�~N����� ���b%l9�%�(����:��L����7>fB��vF��<m�Z�)�~�q"�U�#��l�[����$�E�k�� �~���/��?��`4��4^J�H������C:Wݣ�aN����-܃#��	�Za~v�����=��,����Є�Rz��`
���_��E鹚sHa��Iῒx���.�J�K�{j?���PYFS��f-p��˖�X%��Zb��j��0�x�po����姥�	��q���"��Ԇl6�%��ɥ��Ma'��w���f1d�����at�}>�8���4��jn�Q���/ׁF\�?���P��zo��uy$�Hq��p����տ�1��T�����Ƌ��:��3�7�C�'��#t/t��0Q���.ӹm�FUoz�����,(k=J�*�d�;]�o[<YZk������y��$��O�xvZQ�xr��//�U=M�77 ��$3��/����C����7��Xto��\�i�#x�XJ����$RAN(5䅗���@W9֢o,8I����R�#�	���
AF��0<�0y�J�����`�e��й}6�B�~O��F�??����4Z� �ƭ'''��E���# !H\�c������L�fȁ%,�s���D�F������!k�ڣi�
7S�k�L�r�t}��Ѵ��N��@���d����:�̷��c���U/��9�wIݏ�@�[�����J�:�����-������N�����<W���{�����3�S��'� 0�w�����u5�a�szF��
aǊR�+-O J<�P^%L��5@d�|h.�F� �B�j�߽FJ��5��+�]D��,�i��\)N ��hY��]����&O�����؏�M��G1i�Jm�9sc��s*U���	���,�r�&�T_�P��uI�sV��>q���|l�:�]Q�� ,#gY���@��H{��>p`��	+B�3�:�_)}�@���?]�
�N��gx�OP�p�o��8���uOq�~Ϙ��'^��ƲB�����k{�� ��ܒ\������
��q�>\�b�Rֆ�)������8S�����ny>Iվ$'�c=sgS�t�*_�nGA��-�T,���a���y�ia6�H�j8pv�0\ ذm��5G?~{U�P�&O����*/H��P�eN�7g�����AM��UL@4�����T��~���e����gLr6�*����ڼ��7��##�^W~JJv����я�����:m��@;|n���e+�-���R�s���u'���	�V ���+�R횆&ԙG�7E���@����:UD�h.�.�U��u%��u��T1�nO	«�@ݶ�miɶp��AE K#m��Lۂ�_9$$&��Fvac��h����`K���HW���-���[a�#� ��:��O�1+��)p��ޥ�iН�B#a=�'�_և#kJ�����0T��1�GP��O��r��heKK��H���EKܽƩ�������"^���O��P"�Z+:�G.E��X.U��c��h_i*T�t�ۆ���	�w��d�>�ˡoy���Wz���a+AY� ���zm��B�����@�5�u>�;�K����~��>�����W¢
{�7���*�N���"�?���	�jHt!��3FlЯQ�bԜ��_�#8,��ڒ2��Q��T���S!oe�p�=}3K�/(	���������s�����84aq��c���W���KZZqN���R0�zT9�벗����o�
��Lx����N�es��0/�a��H��T��u�Ww�M)D�z2ۈp�t�R_����ut>]1��	�]���x���:@ٞ��Y+��v���֞E8���T�쩇��RZ�>t�xG�@I�!2��2�i��� �T��	��5�����*vŧ���lR�����_�ׇL����&��	��!F_����b�����j��x�3w���EO��V1F�j�S�Z���7n�(�Z!�D�ywQ)lAs�2�8�yd��W�㠵u�	��V� �K���ؠ�hz�>؁q����y��r����ͭ'�^�����g׌�_eݏ謻bȰ.p{�NrK>��>�Up�~����H�n��
���`��x	GN��A����=���MF�<�����*lIq.�
�E�¯β+�
�N�
�U\|hδ��n!���X��A�����MKGpS^����a��W�Ix������k1� =}��N+�A���1��ZvK9r�t�z�9Z�Z�5�}���)}:`�1�Ϲ�ynu$�k3�(_Mp�1�7���A���
�ow���HX���T��
I3��S����n�KI����?��I�u��S�j u�a�:�Go�_bX�Ù2#�c�L5]R3��6�+i�� �۸}��d6~%C�_���6�7���"���$E鵣Rlׂ�_T���e���VI�!�L.��-i�R�T�E�:��vzn>���*%���k�	�L��a���S�ߜ����]@��?�q���!2�Z����:�����k��p�2]py�4矌E�]�#����g���w����&�2�)��� �㑩����Hjծ�
l!i(	>��i�B*<ٜ/e����c�����L&7�� �������v��GE�PįD��ې��P���&S"SNV�T�5�C��+Ο?p��]x�K ��v\MA�\��7�n.A���0�zG�IC��t�N����i����>�o �4�G��f�RW]��̺њ�?ȱ:]�P�|��#��}c��"��`�U��"]zq���gU�$H݌�ᗷw��:�o �s�0����C@q:@q{a����$�$���O�:��G�cG�� O~���F���s_@waN���s����K�q)��b��N�K6hh̓)}���d�5��������9��+d�lt0���ѿh����__���X��%���c��yhUL�TL����!xᾬ��"���D��-���U�:�U�Y � /��|�ε��0���s�־xQ�Uu6�=��d� m��$�٢mfț��p��ij"W�����i��3Q3��5[���#ȼ��fleW�͔ ��G^�O	���#2]��+3�VI�|�<����;�����t:��(����,��6�L3"s�j�y\�vR�*KKZ�����g;�r�J����BU�Q��:+t�Xʮl��y��}�y���"UġC�L�d��E��#ҏz�6Z�g�����|��+��2q&.�Q� G�8č(poq6�%&�����!l��[�^�)D�!����ǀ�����s^sV�����P�?��:�w�?u��w3�G�v�g��g��>�ڬ��K���c)��<x��2�R{���>�}���]�����<ty,H$�^�K�5E��(�O��:��]G׹�sl&%F�2��dNh�3nXN'�����>|�K7��IDf�+���@s~*=��ت���(�F�5����m�k����ܐ�"��JK[gEq2b�	�W|;55�'s�[�0[mf|@�G^�1J_[�c`�aii�7En���J�XMH5b�
^� .�)2��z	���Y<Q��1Q�$�CS�Sm�p���/��@�(D��ʹ}j~f�Y��䃏��"�CX^�Ծ��y�'�z���$*>��O=tt���Z(U�C��s�aj�\���4a�v%���~l�M��#��9���ĨS��^r�U��o#3pQ�_P�t�R̈�u/Q؅��ܱ����X��<yc����:S���G:�ό��q@1��g���#�Z�Pw;n��7=�O�aA�ߨڒ��02D7�ā�-�5�:�X��vs�>��7N����5�"W�|/�A���"O�����2��	P� X���0���*�x��,~�(P�"��{Py]xF��#�9�,����j@�����j�G�o1��H���?f�W���C�8���wp!1����dv�䩇�t�w���F���y��4�G�����3�>����!k�����p��,m5`�v��ֽ��u%�vq�l��-���*o{qO���+��!zGM�d���9t;'��Eq���`�O�9�$fR�?�F�u�_�N�f�]0�;f��>� 
���x��)x���҉��:+h��d����m6�?��e�m_�&�����N��3�0��R���.]j��&����eSw9B6�������~cV_*,y�g���ǖ2fs�{Vd����n.����B����
�ܐF+�O�R ��������r}RQQQ@#�,Ȥm�����\jj�Y-_hQ����݌Z�h8�@k���0w��.���7��=�Z_dA�ŗ+������"�/MjYa��;��x�xkmo�~ b�pp/�5	�f㣴Ɉ��0���:tmqv�����1��0��h&(-&%�����|�
�����d�'i�c���r=)��F�ϛw}1��ʆ���w�9�ȧ�52�\D�۷,8�[s��r��N�t�*�[�����آ�^hq��g�:Ue���q�$�ׂ�̱�B�Nq�&�ԍ���m��K��R�����q�B��2Bn��(��~7E��Ǿ^;H�#9��5��� �!�����G,�o 2�C�Mք�t�� -�P�YX�'pst2!���HXf�H�2��BZ��:��J�y&z�	D�C��a�v��wԪ���("i���}_�3@y�!Z��U��}Y©�3ؼ;�ݹb��@��O�Hl�P35��;�uB{�.8��k�����%9�zn��)��;Kkǭx�}��d�ڤ���i��+ԯT����'Z՞�N�S�U�'хQ�q�wbƤ���^���w�2��u��ՂO��/����7� �>h�H��}Լ
����!�Iۆ�X�IŢte�	���Cǜͼ�;((�t���f,JeG�eg��z�ѳ�4'2�<t�t�)�b���y�^���9֯�1dM��k�����;Od�#��;�r�F�K�	Up8/�n"-'�kdzs��࠳���:A�����/�0�#h�O>' yn���_1B?UU(&��(��>v<�::�d�^4�1���#\J���Qɼh�?]SC��+��a6������2��6lHh��eY��Jc&��~�ĤLIQf�J���fO����U�ͥ�z��>�c�����]�ni��D��1�[�$CÊ<�g��N������	�}���nb�~j�RQl��j�Ym���g�D:'�W�_GP�5��*\��r�XDۖ��V ����ZnZ�S-Ǘ_�BQ&��D�n���ѣG�����hM��1Q�$ra�!ɘ�L�<m���Uy�S�8��L�Jc�`�R`qϡë_a?��q�#�e�-į��;V��J�8c�ApyL���}�s��=�����T���K�AF��T��o��,B�c���:��/�6A�v�	���y�A�=~|Bq�@B�Z���<4!+"��7sni�{F���|K.L��!2W�qFd��ʹ�t���V�B����<�ˎ[K�����a{�?ǁ�ި�Q!*j��]�<Td������-uw�`P�c���v�����gg�����})9������m�@.�����4��*B��%XEp@��� ���S�� 9X��a]����{XQ&���E.ǢߩcQ�#������Ӿ��^��n\��♰��P���%l޼Y��0��Y�F0���Y��qk�b�k�[�^9j�@G-ѽ�e��YA/Qŧ��}D,^�x��܏�dkFj���>��s���F�"�ᔂ?]5��0��Y;���1�$�1��VO��M�qrs�́XB`�C�PtS���"����,Q�J%�y���ϫ:z?ۗ|��\�~��I�WM��R���x�%0�C�)m����8�/Ļ�&_����A*����+UGC���YS\!b�xV�<'��c��Cɑ��16kn8�9�W	>�O��{��6�1_���4��%���;�W�d�KVڦh`��Aw���Ͷ���M��k������b��7JDG�w��nCOF��n��F^Tc> *8&�+�6�~Z305#�<���#�M|v�cG���#j������F�K�ڡDG��� �R,dq[�T��{M��kY�X��gi#��=�ZRd�C�
����8��K">�� uW�� PJ�}�s����5�R��B���R��l���D�:��W �c��/AK�ɓL	l�!��!T�x�s��ߞ����Ƭ'D�a�5n���5!�9�H��Z+Jj���]��{NKH��0���G:L�}����b�`�3���Yv�B�v�M�O�/I5a� Mi,�u2?7S@�>�^�Ss3�0|
�}�g�$�&f�b%C��t0['6���+���72���R�J�f�����+,�/�  ��d�Z--��J���oI����]��x��)w���l�0F�xE�_y�ou�h�N@��< X*o����k�9Ŗ�"��5��h� �8��ߡkT��S���G7���[M�+������E����#o7P��3I�������� Z����we����+�~f���z��^�Ύ�iALX!�z�Df���g��)�����x94�c�6U}t՗��8��G�*�ɔ���'c�.A�7]Ó�>�(�_)_!k[�ޚ�3�'�$�����`-n�Ӡr�B�-�`m�$?����}�60p5��7�OK��!`*$�g�w�gW|ς�P[�O|�������^����]��˧�r�!����w_�*��X����!��7�抝�Xw����1oZ��;��+�ě��;HX��w˯Y?���Ժ�xqz9OVC=��n��~ۆ�������acI�Ky�5��i�'ȓ_`;�r1���CuJ���O�����_�?#-����2A����XKپ�����N3���g�ۼn����� -�T�����h7�ZR4iK�D� &qqq�(�AǓ�)&Z|��ӆ���>�Q1�����xG�:�Re�~�e�3��8+��W�L�q`Mh++iv��p@ŦM���v���u?&?g͙��L��&_�e��ʛ�Hq^)�V�B��s�z_����l�`s������\�Eb�C���3&=���M5���~S�xn/wl��0r��>>';#o$9Hx��f�=��z��Ǉ�x�`��`Q
�U�2u�^ץ�i�?��0�`?ڡL(��K�� ]�=>_������b,Gp�N$�y5���d����J]��Xs�.���*�ȇ$��Ǻ�٨����z�!-)Vp�ӶN@��:B��fٖ���-/T�̲�q,h�D�"+���{�����?�&Ѱ3� ��ƶ�-���'5�(�H`�*���� dNE�w����C͕+Wdci��63�(	C{�ÿ�5G�pHT��4�:"�2�?C�IM|Ǫ����Gl6�+"� A����߿�n�i�U$}��M��lV�s�������`; ��|�H��i�w�
�,�re���#�q���y�lR�!U ���o_PZ�$Q?d�xٓ?�3I�1F.�q��N��=��kI�5q��l��d��uF�hץ�����\�����w�LE˪�oQ�^�
�"%� �,���݉�ͭ�99Y�I.~%~��LDʱB="�Ž���Q�5xj�3��l��Gy�/1As���_�L�e��WG4��;뵥T;��z�U~ ۞>������>~��k����E�N^s������L�7ջ�x��ѽy�'�On�4�]E�:��*���q��)"�҄}�B�  �+L5J�V����	��0�ӧ�=����+3�o��ֿ�0܍���2���?a�M��h��f���c�e�:f#�b#i|�׶�{A��O]Q� ��F�������fd��B>�Ȭ�"-��.���lMKZ�=9S»!�%�y���h�(&���T
��F24G�����������S���<��z��*%����v��'�	��ؽe�昣�7g���7�a�E�]����۷Oyaq��wϞ=+�T;�l*[!�b0�GF�~_�4u��IF���
�w�>�H�U<�1b%��՘Co�KL��n��S�k����ׯ_G#��&������א�OT�4�u6�̕�n��9�6�����kA�_8��>ĸ.�����}��]u2[���S���I@���߳�@_��##�}Nj��t�Z/��(���1�<@�UU�蜼�:pḮ�K����m��q#6^�df��! ]@'|C$���ŧ6l:�Fzt�7�>گ��j&1���RtQ�V�%E
U ��G�0��$ �_~�҇��9jC(�w�5�uG�����ESx<2Y�P����L�mfc��|���	F|�[���f�:��W�W�v�i�3��{DZY����_��!���b�nĩl�8[G8u�)9Hd���$|�X_Ld��5�w��e�z�g��':c_`�א�8h(m\k{\���B���� ���O/�t�����uՏ�)a� �re�tG�)ҏ��*L���/�䉕j��uDTk�P��A�U�F%	Z�,ɳk�w��7�*�g�٬�y�FVlS�;KZÏp��T3�`G�b�M�� 5�`�z���㧆��*�Dv�VR|J<�0oko�{��ix����\�pd�SK�Oy ���IJ�v���fh^�Ax�7G�l�E	���m�(~�D�9�1�O����q�&'�y~?y����]�o1�/�9\��{m���X/�����
o%��똾��ܐ@��b��%��)k;-pa;�d����MMF���x彏\�7,Ϟu��?Ocb���k;��C�߳���r�/&\�%��js���J���ǝ�<4Dz���Uv��`�[���C�� �C�w�� f�������3��[w��T������	?�E,K���}u�)�ba�6��kTˑ����6�̅�5y�K�	o�c��敿��g�,,+|��/����(�7}O���T�{AH��0:��jjj�J�|���[17���3��xVt��e�����&{Y�#��P��Ç;���5y��݌��<W.�h����Z<
ߝ�+���r��|��Go޼��xaZϑ�bhK�5�3�u�N������=|f`3���͙u��K���#~��y�6#+������,�H�^� ,j����l��������L��F��)��ź�������c=����*rm[*7�,(kA#(�QU�w/�8(���@s��5��Kz��f�'`���y�����%Q�HgNZ�G�t���\��1K�O�+E����~?t~�Z�E�󘻇T� D�A�a6���Q:��=��7�P��CKQ3�f�&5��Gv�{A�C��F���8W��dfb�"O�g��dh�Px�&�_p�fI��(�K������OΘ�K�L�>�S����b;p3Bw�'1�Z�(�)n�p�M�A�/;��(k.�{�3�=g:����V���5���Th�HS��IG��GoN�3R*��-u��݋�I�p�=:��l��{��w�o)9�˙zE�Bz�ҟ���q��{���<z*����2�`�'[�'�K����0�A,g��u�N��T���ۻ�0�B�c�\w?4�R�/�Lߚ�y67����]D�Oh3o]뽕С���3�^g[��_/��������?�a�� �{ʊ��w&O�*j >8���K��N�S��K��)F@����7v�0�߼�ڎ��^�ۗ�wB��y?P�=��/N��ƱMO+��9��A�~#�Q�<�ECA�e.�2ؕ3E��c��G��)+���I�7g<�15iI�� ѧ��Ҩy
�l����Ѓ���"��m�C%�F�������ܼ<×ݺ�n���aA�0����^v�U���r���o�2֋n��84~0�կ�J��wc��r�'ڶ\0���#��NT�����lF+�H�7T/���15a<&�Zߒ�f6V �1_��+R�˷�HA�����4$2�̝��VV]x�
�>G+D��G[@'��m!��ǂ沵���W�Mܹ����.�Y�<�7g3\yPy{Oz�<E䗱����>D�R�Nt�O��3�S���O��&1�A�ɳU��4 ߭$�ALv, ���`bĮ9mM'�NI���V����'�9�xsTn0��Q�^�_F�<(3-�j��ߛq��Z?&���)[�j'��4�	����رG>tγI��#��ު�����r`8*\�b�RB�al.IN�s3T�ο#x���M���vr�ɴ���ݰv��������No���	��_�/�{G�ME�,�����t-f�������5��k�k�ޞ�o!���)ATj����iu�f�ծU��Dr�ģ��Y��B���,��������cmj�K�f��.�z<q��yݒvK�����.��uVRd1���8��q#l�R�6�3u����v*{������D�;.9wUWk*�ם�w̰UlH�Jf��?�&~'�v
��+(�[U�CO���7 �e����7C\�zdlܨ�hN���N2p �Qi�юD�i&GFN&��[XV�KA����#m�@�[
�*�h�h�ͪ��%-��(:�� x���](/ΊX��ď�E��J�'_�z)k>;yb���A��q0���s��
J{��$�l/'AOs�*�Ѩ��2���͙� �E���K���6���8���$&@�U��=70�S&��ޘ��!]6��g����q{k�B����u=��\,�w%~���ܵ��^lS�/=�PuOm���v����=����{n��
&�ށ;�.����-�3�W	�zH��Ĳ������^ւ��"�IV�ָ�7k��$Mp�(�xlj}x!�m�*���Ϟ���YK��vZ�)�GWWWk~@�5����C�?���@��Fj��6o߹�PSC��PUY�B.y��T��0q��l��7�5U�,*������n�ag�&�!��������m�Ő���8����֪ܼ~=Ѝ\�6�<)N�^OWծ�-���cX���#U/�R�c�+�D�G��\����T�:sj'q�I x-��$��=�TWW�l��X��|S8,j'Dc#"�1L}l����I/$�<�Ƃw:H`����
O��9�sZ��<��r[���q��i�\���x��-ĳ}bi��?Ԃ�}?�Nv ,��CE_T�M@LJ��`�%��MH�޲+��ߢ�Q~�
T7L�9Z��xq>n@fLd�����֓���e<�,�Sq�U������K`�Vv܅ͼ��5�Qmy�����B!:@�v��i�� �%�W�x�Xj�v���*r�0b=�����ק��t6n��'��/�pB`Js�1z�mqU;�.+��rZZ���\ɭ��4���%�~�HC�=\���l��r����x��%�v�S��p�G��=��Jb� �S�e�'��~H�8�֎.i'��_q"�d�����F��=�S˹l��ޑ����Q�����4a'��r��cݫN���z"�B���.�o��+�c���7��<�ס�?,�8�Փ�C8��K�� �Q��c$9�&^K#���	,'�g;�[�(��V���EShim�������-�)46���sa��vf��)D�#I��u$���$�~	�t3�V�K^��b�LD��Wp�L��*���S*�\�~���dp�v0-��4��� �\~;0nҥ�P�F���
�[�n%�s�B�T	�.	,�7����fM�a"7d��W 1z!Ъ�W?t�)�&����玠�|�}���ld�!��3p� �#O��:��.9X__o�@����<Y�a�+��3�Y|�1�旧�!���[
p�R����Ƶy`�/�}~vA��D��6���z�33v�^wez��Y�5wLsQ'.[R�>�7W,�����$ܡKz���)�s4~%��-S�L&S��[מ�lm=R���ڶ�]�y�H-���S���K�@����\�.��@7���-В���m,U�e�������e-K�l�2�o{!�I�ٳg���z���z�	��T;޴X��wU��04��;�I~�����*M���*�Q:�ֵ� I�e��ھ1v9��a?ul�8kn�a�m��DZ�!�u�y#�WgC�¾(��,88�̛>��Gq���K�D��c�)q�ϢйN���7y�a/��o11��1� ��D%t;�m������p}7+�	%=������,�ʛ����<����t<����.�sr���T�fG�t�P&č3�����I,|����Y
6��І�5�ǔ��N'Q N���#Ʋ+U�Fy@1�f�}u�wѫ���]U)���X�MnIE�
Z[�c�/�k��闬����ݻw#cD���@�Z~婭�!;��Ű�r{j�t��Al����r,��16@7$�����7q�;�
\�/��Ѭ�H�.y{��E@g�G�M�X�겗����t@����0���p�1,�w�k/�b�vv�
9B6.�GbIލ�U��F����$�J�D��b��Ɂy�&ѧ�rN3�'Ķ|عUײ�D�������@q������)�ě�A�S}KZ͆^p�A ����7��1�o@�.l���,9�Rߗ1\�*�z9�ߡ+��q��(/,�d�&�(Kc�������g,�-��n�w�F��|���3���؊c��5�_��q��k틆�¤��C`&:�������5�����*�$��s�Z�x��BO�wɛ�,�*��]�>���[N�gk���UV߷ۘ�X��ly.~�H��Y,[�u~�:����ٮ�!-]?�Ə�|9��9�)���y�5�&�F�kO�|�2������酱�Xg������Nz��ʔ�Tl&t� ~�0��X&���xs�����nB��vY��O�0��U�����8�猫>�Ϡ�ȓ�Ad�w�~k<KE��Hd��%_������-���N��.j�kk�e��V�[qz�NB>�1�Mx���DIY��=He۟-�rj�2���7A#�D!\<J�v�p�'OD���C
$��{O८���2�%��7M"�.[�n�h��V�z��c���Yb�	x�?h��H���a�%�L���m��NjR0_��P�E!L'���\�,^��A�cOI�(>H�
�8��aMg�ys,�>����~;n�p�9��H�=Ԇ�^�A�!�9�G����� ��P�՞��@I^J���lgpx��C��8*��	Y��C�R,�a�?~�x �4�{d �����,��;k{��]�2t�Ba�n�h���Yj�J���4s�W�"�ը�guX���	+*cU"\u�r΂n%��J��/�0����_����F���_��w����u�I����i�v�A�܇+���b�m/��[�X��1[����YL�[5sQ��PMu~*��sR�mf�M1�Ď5����큘a���� ���@��zU���p����
s:�m��';�f�lN�����i-@;y;�B`����]�fo#+�J%C�Y��iac���+����K�bͬL�P�_��o)!2S���b���6�B���`ᄛ7g��'�s(�5�{4�_�H	����3�a@;8S[�ݴ/��+ �&�l���I��t�F������{D�/-��^ԛa�-[�� !�R�Ap�ͦ-�9n���2؅�Z2[���xT�_�x�hA���3o�l� kS}spPrb�>d��j�}]�x�?�KΠ�^�����G��%&������
��!�U��s!5�y~�j8�,=�qi���'0H*y{N��uܛ�P�߾v�AAqVvi�x�:[�&������مm�"r�g3gۑ|��k�[R��|}C�,�lb��9�qP��u3�Z<���t�%�"�����\��/ֈ=H�FP���-^�3)V�f�
	��צD;{8D9��V�@���E�ü�ʰ�պls��d�a�ϙAP�4D���7'��n�KǼUH�R�e0��k�gmQٴ��5-��Ӷy,߂i=*/��S�yj�"Yhz�r �>����:�0����Nb(�5y��OR���d��*�b7�P�6�Q�����C!��
���7ޒ��w�| �C�z8��ա	��������A��,�R3K����.�,;��;��-H�u��=�I�5k�4� d �ȱݢ���/��ЋJ-��\���j?Wqnx��˒Ƚ��(��=S��{ �މ>X3�)�dE5ʡ�v.��Y���Va�جP�;��Cf{ O���̲A�G��h�Bn��=mf -�>R��䰊����$��C��]��X����@��w;;���՗`-굫I<'�w�\�w��})�l��	l����S��,�J�ld�քJ�%���#����1��,��:�eb���f�	ÕH�{��ڂR���SCհE�%�eb���3�>���ϑ��FLHC��l���é���!&%,T����#RҬ����%�->���"��֪�oaֱ�>=��ehG�ai�2��v[C֒`=�̂D��K�ڃm=!g��ܛ[��a�q�W�K�1�<)�� ;��o4#ZA@�ӈ4�Nt�.�T 5���v7�Z~�n_��8��ff'U��޽{w�||�C�%=M�Os�=WY�Q �;��p��*ȐëH�U��}�&�e0���ŭ��Wܡz���R��X�[*�^�����m:�r��G��yM 
"MI<too��/|�Yb�^'+��&�ƛ]�gu�b�7����2P�}��r��p�T�ٗ!��VRZj������w�d���$[՘�us�~����X?0��^���/����7nd���ev{}W�D��*�"�'X�B�F�r��kf���z�D�b��k�Gw���gv9|�q81��`f��h��h
E;���K������N:�VUU5#S!�MwƤ�e	*	��[���t3 �C�iB�Sv��;��)帾�1Q`�){U�5�ւ��3�`�,�;tsO�7K1�~K�GI���D�8[�����tU���Y�c��%�*�<F��$	�!��l-�;'BA�����܈�F"����#|�c�h#��ݴ���l,��pћ������=����7�Yr�..��qէO�\�:Q1�c�7�}!�}�q�  ���}&�yP���Q�ekU��'�`��)�,1J�ꤢM���#9�F��y4�:��lKk��z`{�]Ix�XwYkmml���CQ�9�a�Ო2K"�l.����:1��Z��T��1��SCʅ*�<uUS�ec�����t�3���!?�{�n�G|f2����ě�_t^]��gW��fT��)����U�R�XJ���c��f��V�2`D[�w��P�� G(�v�l�K%���Y�1�6
�t�'-.v�?Y�v
�=�uߛP�S�?\By���C���~̦�d��G��e�5�G�W|ڂx�鴦�s_��K⥣��?	��Z�4h �a���|�}�>���<9$�zc6�=d������j%������%���P[kfZ?S���Q�?��Jh��,��[���|�I�rh�Ɓ�Ȅ����Y�tD-pf��\~�6��MnC޲��X����2/��:���rzO�?���D����;�/~8�c�޷���B.o)���(���������}�8�I)��底*�������q���R/,��������+�/fC��:��s؋�Ʒw-�O$�T�4��h.,��iyY�яkzū1rb�bxI���WzX�UG����@nl/�w�kM�X/��y�6tͲ�?0�p�W��n�_�^�⌸����E�FK"�v���\�6ydggW�닂�#AZ�)1�ֶ�kl������X_e'F̷-����M7�)D�!����ٗv�X�G^�ûV��Dol2Q7gf��;��`+ۘQ!�~D�o��6I�]��=��g����0[냙y���*k��g�m\�+�ޙC3N~5��6�r?�O�us���bۼ:Ͽ���o<��t�n֧T����a9����E���X]]}���z*Q������I7�������Q1��$v'�1n�Sq��l[☝�X��-v�w�[o(ě����I�L@n�����
U��Nu����Ʒj�')�/��z.�v��(���R6��gۖ�:����e�c�k���̓&C��S�gD��e:�R�yS�d���aas��b)�Ĵ]���مY���vT佰,��'O�4N�k���:U�����^�����y�<�rN���؇������{��1�M"2L"�ah���+��"g�)HK��-/�\@0ܧ ����-�UG?U�R ���ߦ���������S�~A��	÷���YlX�k�˨$�2�lT����~��s[hZ޸/ҟS�MΙs���?�)�J��F?_�m���14�O���$��/��J4�͵r�{����9�7==��2^O ��rm�°G�`�y�o��b�+7n�:a�9�Ӳ�z^��L�C̢�>,�<U���=�z���o�d�+���YVo�S�6��|}�6y���Z��ktnX>O�%�n3;��8m�׸rQ��r����(Se`/����~ �a�R�"�
���n[>?�����O�<�v�^�hu���Ѿz��`8�Sj ��mll�O}��IY|e"s7(��(ϋG m��?[��ڧO�Vg橋iy��V*YG����z�`/�`�:������կ��)~�a�g�kl3�#e��+&�5�?�{]���4��T����5i=��{4�����@p���2������%=�Ez��g�c�]4��ٍ�Ѡ��e��)co�R���-�~X��C��;�:7F'�E�׹�/#o���n�l�ZԞgG\]�VLz �z�pի�_�v�$�9cb�f�C�LF��p�2�����ބUS�866�K���"�2x�4�~�i�ymch�zrQ�Ϝ�W��k䐇�[hA��5<�&�����z�qi���pܢD����̤/��9��?k���%ej�n�
��h��bQ�gm\e�_h}S�2����&]FeD�?5�����?��i�����+h�o7�`�<��W��V�`\��.X �Oo�Mzۗ�
h���E@���;00�N!� R���gU�puum����T�����4��0z�OC��z���o)a˻��S��1zy:U�Nm��!�.Z�hmk@����3hJ�hJ�����
|H̑��^�f������-�Bw�g?+J���C��VxY+�;���#٨�WQ9��j�'B�ҽ5л���$�*�%Y���cJ�D*��$��u@�o�Yi�)�|�Qa���,��b����&�*�,�Sm���EC���?bE�x�����I����@� f�`c.q��9X䲰�ۍo)D���X�h���^������>��ؒ��/�-j�x��5�?X
{Yk�Tq?���k����@K� ������� �k&�tǎ/N��LȞ�| z��p�ݢ�]�L~�;`��k�9��U��?F�z�G��_�J���E=y���4�)�E%蹬�Ud�w09��D�ٴ�&FA//�$��f�%&xA��`�FR��ar�H@;�~�Z�8����l�%���������m��#��
߈�>�yg�e	F~Tﳵ1���mh�ݨ{Vl���WL�s�b�?��%�����o��Y�$��Z���_E�}�G"����o���~v|��.������_����]����u��M�ǿ�+ǰ�tP-��?f�����y��ù���̼f��7Z�m����,��1����_c����]33ή���GI)v��)���?��y~���+m3��Ϡ�:�f˵���^��CZ,�{���0;,{-���p��Mn}��g����f�}�[�zD��l=�/.�:�._��[\GL�ՠS�<jv���-���	�K���^�U�d�ګ���W��\�v$�{B�@y���ӱP�ս��nª6��\��	���%�~݃�D�}ՄA]�踸o��=�b���_�y��ZkZ�ð3'7w/�p�~������ޯ��v�^\��L���a�����
H�j��:-H��Btiv�k�X�TK��+Q�:����7��ޝT�Y����Q��|_̏z-�ݿY>j�@ݠ:���O=H���:���v��� =N����M[�0�;�-<�nݻWWu����ph���zOj�Z�]A^�{�J�!=�/׼ ���ֶ�����\����]�E�z�_��(�S����r�V.pvj�\[�v���O��KB�7��Q�a)��o��2�ʾ�Z���Ũݶ�`��� S�^{]�Z}љ�#�F�k�Fâ�t��RPG>�����Ӡc9����T�_�
JUo�^�)'����_`��Wr���Dff���`��f�����}�]w�Fłba�Z�x'���Ps�^�Ut=
�'=\a�MU,�;_�_.G��/���&�k������)�	 PK   �XXʪ��;  6  /   images/1a471211-da5d-49df-af40-e9b794edd793.png6��PNG

   IHDR   d   �   5��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��pW�	!$�RB���4���H��dG���P���m*�V�tZA������c�H�D�8�V�TfJ�"��B�_����ޣ����{o��ݻ���Nr{{����������Q�5j]�p!����g�g�}={�J�H�Pv)��]�|M����~�}�}�}��&� ��ىToz��)
S��ȑ#/�/� ��5�O�'��ag(_�t{�Z�y��i�?�{�;ٻ؇(	���sɀx��G8���3ط�od���@$�']�~����+{3{#{7��B��u i@\Ǿ�=��A
W%�%�Mv3{-{�_b'�=�&k@Ҁ��~�}��uSҀ��]On��(�`�$�	�`�F�:�$̳�?�'��%P )@�W��~����@��Y��o���و��������4{��٘O.�%��AFK @$W�W��Snj4�g������7	 �fWP�����V�o`CP|�`|��I!叐E�Ʈc��~��`���姐x��(�yl�����Rh7�~AO��6�Ք��!ȕ��&P��H0j�m3�zk5����.�6��ʯ\U���-�8�]���@��X�KV��rG��@'JL"�N��d՟�`�Dn:_YJ@<с�����ı�	�%�r7��S+5�An�{��t�<FV�z��⩮0��I������'U�-�AⰘ�t�3'�z��u�L!+SM���`��Cde�I�;����+��TDc��ߎ�@�謌�Luy���8���[�� R<��RZ�,�@V~��\��cF���H$��X���O�6�ZeY >� ���/�L8n������$�*K@��.����Q:~J�^%VfU)Y�L8v �z��sY޶�J]��tNh���':�gEh̵��"�[�/���'��"%�ҍ�"$���V,��F�[u�N֮�.��A�a���Y`�ý��0LOV�� ����IV�I�;L���ĉ��J
�dذaN�a*ߗ�Y��7;zV��Ȫ�,�����,�����,�����B2t�P***R�`���Ң��2d4H�}Z[[�ܹs�B2o�<���t�*B:����8��>�f͢��j��+`8�֬YC;w*_��B�����L��e�uM�����尪�%��'�W��\*U��U/b�F��
;d�����b�d�@� ho�M�F'N�ո�>y�$mݺ�rA��ƶ���O�n*��HJUe!rr�*��|�1�<�D���s��Ç�y2��b{ 8�cƌ��K��|��85��a\�D%䍆8^��@�T������ �"$b�4Щ�E��S.(6@�po۶��?�kF+����iʔܸ�]l� 2v��E����S�Nu�O�|�wl�@���mϕ��
H>���r�X&�m��� �N�>�g;@<8V	Ɯ r��є�E�M�Ν�\��8%'� ���ё�]K�@2� f]�7Y Sh@0�F�GeE��֚T?��ŊvUa_�U�A)4 [�l�ݻw+��		�����8r���:t��Rh@���.���ݻ�q\�
$��hK��I7�J$G���[^z�~MJ���_�@�+3n*֦����O�����D�e�U�Qȿ�1~=���
u�����]+}�R�Q�M���de�ߪ�d�?��b����*#���u�����$�5�<��~�۹uk6~-�9��d$LU�t^�����=��T�<�-$EU���SmAO�g���U&e/�?�f�9sF�E&#o�B��^IV��5r�oZR"E��ٵ�;�&��������Jc.�!^(���s;::v�_�HX&B|,�())Y(]������ﰺ��g�0F�=���UUUO2$�r��kپ}����v$�2M�u��������sw�cǎ5�ٳ��Lӆ=#F�(���~���Pyz����mǎ�[[[[������k�ٳg�0j"m "J���p]�~���q�&M�D+V��j߾}5�mݴiӲq��ubf/��O�N3g�� '�|^>0�oذ��7oN�τ	��������q�NV[cc�����Ç;��x �nt@F"�8qoB�9s�Psss�Aq�t����-J����˝�E���g��ŵ���	H]]q�����೗͟?��'&�	�['֟��F�d�DL� U
�g���8�\!��f݋x
��}��o �耞���z�N<�(�D���}�A1����o�+���9�4_7���~�B1"�@
�4�u�WddYX��9�a�E�k��~��`��^G�p�@�"��7x���_�o'w����A���B�MH�cF�d@(����_��`��
���w��&P���p	��U�o�p;۹�}D�h��o4|=� ���F�sܐJY�d�RJ@�*
�|�R��/^La	gq�;�a����←�ȋa�۹$B5Z�"���?&7:���-=��}/�큩����*���P����L�|��?�x�ׯ<Q�g�z�
��~�=���l�/��%-	����M�_X#|)�uIo�`o"��g|����SrD�	J�7�`L$w=�5�_Xz�^L�������u��ȭZ�
��½��+�P� �`Ԑ�[b�"�)��F�!J0�$(��m�@�8��h�w�RA�D�����d6r��� �ubCaIP�����P���vd����E �*
F;����bC�aIP�c���	e��W�r�&��q���R$6xt�mF0����!6���m	�]�`�Y4z^h
>�v.-P�6^!��=�M����CH���VrS,�}���dy��ERt �a�/D�lJ҇�CH��<է�����B9(s*�{x#�,�ɿ^fב��8���������Z�E#ł��ic��wɿ����wC.����=Ay�{|�BqAT� �${T ����!	
�~t��|�G���� t%� :$��!	
�(u�v��Q��U �	�+|��˯z7�2!	
�+��K�˰H��n�>>�G�����11�;�G��@&���%?���o��`a/RD���o��!�ko{?X�J��)`̃�2(�@L���3���@�.	��)5���N�<�� V�<P�����@����>��O{ȝ��� �I�FG
y��� ) {���^�1Y �1���B\Ez�Y�U`ڨ�w/n}�P|t��~xI�B�    IEND�B`�PK   �XX$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �XXP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �XX.�&�  �     jsons/user_defined.jsonŗkk�8��J�]�����o���f���.e�e�58v�KK)��{l��Nme30�Yzt,�=�/A��"hk[}Kl�6	f����,���9������u������Zo���*i��<�^��D�{WV�01����4e�Te��*����v�,R��vd�3�,��I!0��1�Q3�BrN�q�lm�l�A���3�SN��1#�	Q(�DR��N��r�-�`]�w=��B?V��(��6+N��/A�nVY����q��]�j.`�~��|��ɰp8���Z��8M.�*���8�	e�u��r!L��݃�^澬`I�h��&ױ�f]��/OV��lK�X>��������K�Xᅽ��m�X6Ɔ^X6g7N*S�U��b̌����+C�OC�J���\�h�^�%v2՘�P�G&q_������_R7t,*�w���K����%wCǂ�~W)�б���3��<��N(
{bWK7vBS��<� �XV��q����E�vE\����ź�@'���źEK'�V�u�:Q��'V��5+�Fn�Xc}���J7u�1J<���:�X_|��,C'��"�(\ܓ��(]�V��]�'�-.6Q��'�u۷�W�7x�*h�_a��C�mB�Qd"�gQ�b�л�)��$���{[�[[5��:��F=
=��!6ۢ�:o{GQⰻp�nͮ��/�Ί�r�}���7Y�Ź}��C���7���v�E�jӴ��m=�_�5���%ea����O8ō��_J�I�y��g��hso�����Z����*]�Yݔ��ǟN���>�>�!o���ƈ�Ǆ!͒a��b��XY_o�����E� nc���q���K�}�����)�]5�j�\)�xP<�[[$�9H�ymtt�G�Έ8ɃVj*�I�QE�y����b]ۃ�k"
��S&�P(�I���M�4�����*�M�^0e��A�SƦ|ԝ4�KDsI(!(�`͹JR�S��U�T�&�T�'��?WC��9c�����N3�]y���?PK
   �XX��$x�  �                  cirkitFile.jsonPK
   �XX��8��9 z /             '  images/07769342-c5fd-4eb7-a5a5-41db20f507eb.pngPK
   �XXʪ��;  6  /             'M images/1a471211-da5d-49df-af40-e9b794edd793.pngPK
   �XX$7h�!  �!  /             �Z images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �XXP��/�  ǽ  /             �| images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �XX.�&�  �               D/ jsons/user_defined.jsonPK      �  |3   